  reg [15:0] q0, q1, q2, q3;
  always @(posedge clk)
    case (a)
	// foodfight code 136020-302.9c, 136020-301.8c
	13'h0000: q0 = 16'h0001; // 0x0000
	13'h0001: q0 = 16'h7578; // 0x0002
	13'h0002: q0 = 16'h0000; // 0x0004
	13'h0003: q0 = 16'h008c; // 0x0006
	13'h0004: q0 = 16'h0000; // 0x0008
	13'h0005: q0 = 16'h008c; // 0x000a
	13'h0006: q0 = 16'h0000; // 0x000c
	13'h0007: q0 = 16'h008c; // 0x000e
	13'h0008: q0 = 16'h0000; // 0x0010
	13'h0009: q0 = 16'h008c; // 0x0012
	13'h000a: q0 = 16'h0000; // 0x0014
	13'h000b: q0 = 16'h008c; // 0x0016
	13'h000c: q0 = 16'h0000; // 0x0018
	13'h000d: q0 = 16'h008c; // 0x001a
	13'h000e: q0 = 16'h0000; // 0x001c
	13'h000f: q0 = 16'h008c; // 0x001e
	13'h0010: q0 = 16'h0000; // 0x0020
	13'h0011: q0 = 16'h008c; // 0x0022
	13'h0012: q0 = 16'h0000; // 0x0024
	13'h0013: q0 = 16'h008c; // 0x0026
	13'h0014: q0 = 16'h0000; // 0x0028
	13'h0015: q0 = 16'h008c; // 0x002a
	13'h0016: q0 = 16'h0000; // 0x002c
	13'h0017: q0 = 16'h008c; // 0x002e
	13'h0018: q0 = 16'h0000; // 0x0030
	13'h0019: q0 = 16'h008c; // 0x0032
	13'h001a: q0 = 16'h0000; // 0x0034
	13'h001b: q0 = 16'h008c; // 0x0036
	13'h001c: q0 = 16'h0000; // 0x0038
	13'h001d: q0 = 16'h008c; // 0x003a
	13'h001e: q0 = 16'h0000; // 0x003c
	13'h001f: q0 = 16'h008c; // 0x003e
	13'h0020: q0 = 16'h0000; // 0x0040
	13'h0021: q0 = 16'h008c; // 0x0042
	13'h0022: q0 = 16'h0000; // 0x0044
	13'h0023: q0 = 16'h008c; // 0x0046
	13'h0024: q0 = 16'h0000; // 0x0048
	13'h0025: q0 = 16'h008c; // 0x004a
	13'h0026: q0 = 16'h0000; // 0x004c
	13'h0027: q0 = 16'h008c; // 0x004e
	13'h0028: q0 = 16'h0000; // 0x0050
	13'h0029: q0 = 16'h008c; // 0x0052
	13'h002a: q0 = 16'h0000; // 0x0054
	13'h002b: q0 = 16'h008c; // 0x0056
	13'h002c: q0 = 16'h0000; // 0x0058
	13'h002d: q0 = 16'h008c; // 0x005a
	13'h002e: q0 = 16'h0000; // 0x005c
	13'h002f: q0 = 16'h008c; // 0x005e
	13'h0030: q0 = 16'h0000; // 0x0060
	13'h0031: q0 = 16'h008c; // 0x0062
	13'h0032: q0 = 16'h0000; // 0x0064
	13'h0033: q0 = 16'h0112; // 0x0066
	13'h0034: q0 = 16'h0000; // 0x0068
	13'h0035: q0 = 16'h0148; // 0x006a
	13'h0036: q0 = 16'h0000; // 0x006c
	13'h0037: q0 = 16'h0148; // 0x006e
	13'h0038: q0 = 16'h0000; // 0x0070
	13'h0039: q0 = 16'h0148; // 0x0072
	13'h003a: q0 = 16'h0000; // 0x0074
	13'h003b: q0 = 16'h008c; // 0x0076
	13'h003c: q0 = 16'h0000; // 0x0078
	13'h003d: q0 = 16'h008c; // 0x007a
	13'h003e: q0 = 16'h0000; // 0x007c
	13'h003f: q0 = 16'h008c; // 0x007e
	13'h0040: q0 = 16'h0000; // 0x0080
	13'h0041: q0 = 16'h008c; // 0x0082
	13'h0042: q0 = 16'h0000; // 0x0084
	13'h0043: q0 = 16'h008c; // 0x0086
	13'h0044: q0 = 16'h0000; // 0x0088
	13'h0045: q0 = 16'h008c; // 0x008a
	13'h0046: q0 = 16'h46fc; // 0x008c
	13'h0047: q0 = 16'h2700; // 0x008e
	13'h0048: q0 = 16'h207c; // 0x0090
	13'h0049: q0 = 16'h0095; // 0x0092
	13'h004a: q0 = 16'h8000; // 0x0094
	13'h004b: q0 = 16'h3010; // 0x0096
	13'h004c: q0 = 16'h2e79; // 0x0098
	13'h004d: q0 = 16'h0000; // 0x009a
	13'h004e: q0 = 16'h0000; // 0x009c
	13'h004f: q0 = 16'h207c; // 0x009e
	13'h0050: q0 = 16'h0095; // 0x00a0
	13'h0051: q0 = 16'h0000; // 0x00a2
	13'h0052: q0 = 16'h20fc; // 0x00a4
	13'h0053: q0 = 16'h0000; // 0x00a6
	13'h0054: q0 = 16'h0052; // 0x00a8
	13'h0055: q0 = 16'h20bc; // 0x00aa
	13'h0056: q0 = 16'h00ac; // 0x00ac
	13'h0057: q0 = 16'h00ff; // 0x00ae
	13'h0058: q0 = 16'h303c; // 0x00b0
	13'h0059: q0 = 16'h0000; // 0x00b2
	13'h005a: q0 = 16'h207c; // 0x00b4
	13'h005b: q0 = 16'h0094; // 0x00b6
	13'h005c: q0 = 16'h8000; // 0x00b8
	13'h005d: q0 = 16'h3080; // 0x00ba
	13'h005e: q0 = 16'h227c; // 0x00bc
	13'h005f: q0 = 16'h0001; // 0x00be
	13'h0060: q0 = 16'hc040; // 0x00c0
	13'h0061: q0 = 16'h7e2f; // 0x00c2
	13'h0062: q0 = 16'h22fc; // 0x00c4
	13'h0063: q0 = 16'h0000; // 0x00c6
	13'h0064: q0 = 16'h0000; // 0x00c8
	13'h0065: q0 = 16'h51cf; // 0x00ca
	13'h0066: q0 = 16'hfff8; // 0x00cc
	13'h0067: q0 = 16'h4ef9; // 0x00ce
	13'h0068: q0 = 16'h0000; // 0x00d0
	13'h0069: q0 = 16'h04ea; // 0x00d2
	13'h006a: q0 = 16'h303c; // 0x00d4
	13'h006b: q0 = 16'h0000; // 0x00d6
	13'h006c: q0 = 16'h807c; // 0x00d8
	13'h006d: q0 = 16'h0004; // 0x00da
	13'h006e: q0 = 16'h807c; // 0x00dc
	13'h006f: q0 = 16'h0008; // 0x00de
	13'h0070: q0 = 16'h33c0; // 0x00e0
	13'h0071: q0 = 16'h0001; // 0x00e2
	13'h0072: q0 = 16'h861e; // 0x00e4
	13'h0073: q0 = 16'h207c; // 0x00e6
	13'h0074: q0 = 16'h0094; // 0x00e8
	13'h0075: q0 = 16'h8000; // 0x00ea
	13'h0076: q0 = 16'h3080; // 0x00ec
	13'h0077: q0 = 16'h207c; // 0x00ee
	13'h0078: q0 = 16'h0001; // 0x00f0
	13'h0079: q0 = 16'h73e8; // 0x00f2
	13'h007a: q0 = 16'h4e60; // 0x00f4
	13'h007b: q0 = 16'h4eb9; // 0x00f6
	13'h007c: q0 = 16'h0000; // 0x00f8
	13'h007d: q0 = 16'h897a; // 0x00fa
	13'h007e: q0 = 16'h46fc; // 0x00fc
	13'h007f: q0 = 16'h2700; // 0x00fe
	13'h0080: q0 = 16'h2e79; // 0x0100
	13'h0081: q0 = 16'h0000; // 0x0102
	13'h0082: q0 = 16'h0000; // 0x0104
	13'h0083: q0 = 16'h4eb9; // 0x0106
	13'h0084: q0 = 16'h0000; // 0x0108
	13'h0085: q0 = 16'h7bea; // 0x010a
	13'h0086: q0 = 16'h4ef9; // 0x010c
	13'h0087: q0 = 16'h0000; // 0x010e
	13'h0088: q0 = 16'h008c; // 0x0110
	13'h0089: q0 = 16'h2f00; // 0x0112
	13'h008a: q0 = 16'h48e7; // 0x0114
	13'h008b: q0 = 16'h7ffe; // 0x0116
	13'h008c: q0 = 16'h4eb9; // 0x0118
	13'h008d: q0 = 16'h0000; // 0x011a
	13'h008e: q0 = 16'h102a; // 0x011c
	13'h008f: q0 = 16'h4eb9; // 0x011e
	13'h0090: q0 = 16'h0000; // 0x0120
	13'h0091: q0 = 16'h8048; // 0x0122
	13'h0092: q0 = 16'h303c; // 0x0124
	13'h0093: q0 = 16'h0004; // 0x0126
	13'h0094: q0 = 16'h4640; // 0x0128
	13'h0095: q0 = 16'hc079; // 0x012a
	13'h0096: q0 = 16'h0001; // 0x012c
	13'h0097: q0 = 16'h861e; // 0x012e
	13'h0098: q0 = 16'h207c; // 0x0130
	13'h0099: q0 = 16'h0094; // 0x0132
	13'h009a: q0 = 16'h8000; // 0x0134
	13'h009b: q0 = 16'h3080; // 0x0136
	13'h009c: q0 = 16'h3039; // 0x0138
	13'h009d: q0 = 16'h0001; // 0x013a
	13'h009e: q0 = 16'h861e; // 0x013c
	13'h009f: q0 = 16'h3080; // 0x013e
	13'h00a0: q0 = 16'h4cdf; // 0x0140
	13'h00a1: q0 = 16'h7ffe; // 0x0142
	13'h00a2: q0 = 16'h201f; // 0x0144
	13'h00a3: q0 = 16'h4e73; // 0x0146
	13'h00a4: q0 = 16'h48e7; // 0x0148
	13'h00a5: q0 = 16'hfffe; // 0x014a
	13'h00a6: q0 = 16'h207c; // 0x014c
	13'h00a7: q0 = 16'h0001; // 0x014e
	13'h00a8: q0 = 16'h86dc; // 0x0150
	13'h00a9: q0 = 16'h227c; // 0x0152
	13'h00aa: q0 = 16'h0001; // 0x0154
	13'h00ab: q0 = 16'hc040; // 0x0156
	13'h00ac: q0 = 16'h7e2f; // 0x0158
	13'h00ad: q0 = 16'h22d8; // 0x015a
	13'h00ae: q0 = 16'h51cf; // 0x015c
	13'h00af: q0 = 16'hfffc; // 0x015e
	13'h00b0: q0 = 16'h207c; // 0x0160
	13'h00b1: q0 = 16'h0001; // 0x0162
	13'h00b2: q0 = 16'h75e8; // 0x0164
	13'h00b3: q0 = 16'h227c; // 0x0166
	13'h00b4: q0 = 16'h0095; // 0x0168
	13'h00b5: q0 = 16'h0000; // 0x016a
	13'h00b6: q0 = 16'h7e7f; // 0x016c
	13'h00b7: q0 = 16'h22d8; // 0x016e
	13'h00b8: q0 = 16'h51cf; // 0x0170
	13'h00b9: q0 = 16'hfffc; // 0x0172
	13'h00ba: q0 = 16'h4a79; // 0x0174
	13'h00bb: q0 = 16'h0001; // 0x0176
	13'h00bc: q0 = 16'h8a7a; // 0x0178
	13'h00bd: q0 = 16'h671e; // 0x017a
	13'h00be: q0 = 16'h207c; // 0x017c
	13'h00bf: q0 = 16'h0094; // 0x017e
	13'h00c0: q0 = 16'h8000; // 0x0180
	13'h00c1: q0 = 16'h3010; // 0x0182
	13'h00c2: q0 = 16'hc07c; // 0x0184
	13'h00c3: q0 = 16'h0080; // 0x0186
	13'h00c4: q0 = 16'h670a; // 0x0188
	13'h00c5: q0 = 16'h4eb9; // 0x018a
	13'h00c6: q0 = 16'h0000; // 0x018c
	13'h00c7: q0 = 16'h8902; // 0x018e
	13'h00c8: q0 = 16'h6000; // 0x0190
	13'h00c9: q0 = 16'hff6a; // 0x0192
	13'h00ca: q0 = 16'h4eb9; // 0x0194
	13'h00cb: q0 = 16'h0000; // 0x0196
	13'h00cc: q0 = 16'h8048; // 0x0198
	13'h00cd: q0 = 16'h303c; // 0x019a
	13'h00ce: q0 = 16'h0008; // 0x019c
	13'h00cf: q0 = 16'h4640; // 0x019e
	13'h00d0: q0 = 16'hc079; // 0x01a0
	13'h00d1: q0 = 16'h0001; // 0x01a2
	13'h00d2: q0 = 16'h861e; // 0x01a4
	13'h00d3: q0 = 16'h207c; // 0x01a6
	13'h00d4: q0 = 16'h0094; // 0x01a8
	13'h00d5: q0 = 16'h8000; // 0x01aa
	13'h00d6: q0 = 16'h3080; // 0x01ac
	13'h00d7: q0 = 16'h30b9; // 0x01ae
	13'h00d8: q0 = 16'h0001; // 0x01b0
	13'h00d9: q0 = 16'h861e; // 0x01b2
	13'h00da: q0 = 16'h4eb9; // 0x01b4
	13'h00db: q0 = 16'h0000; // 0x01b6
	13'h00dc: q0 = 16'h7468; // 0x01b8
	13'h00dd: q0 = 16'h207c; // 0x01ba
	13'h00de: q0 = 16'h0094; // 0x01bc
	13'h00df: q0 = 16'h8000; // 0x01be
	13'h00e0: q0 = 16'h3010; // 0x01c0
	13'h00e1: q0 = 16'hc07c; // 0x01c2
	13'h00e2: q0 = 16'h0080; // 0x01c4
	13'h00e3: q0 = 16'h670a; // 0x01c6
	13'h00e4: q0 = 16'h46ef; // 0x01c8
	13'h00e5: q0 = 16'h003c; // 0x01ca
	13'h00e6: q0 = 16'h4eb9; // 0x01cc
	13'h00e7: q0 = 16'h0000; // 0x01ce
	13'h00e8: q0 = 16'had94; // 0x01d0
	13'h00e9: q0 = 16'h4cdf; // 0x01d2
	13'h00ea: q0 = 16'h7fff; // 0x01d4
	13'h00eb: q0 = 16'h4e73; // 0x01d6
	13'h00ec: q0 = 16'h46fc; // 0x01d8
	13'h00ed: q0 = 16'h2000; // 0x01da
	13'h00ee: q0 = 16'h4e75; // 0x01dc
	13'h00ef: q0 = 16'h46fc; // 0x01de
	13'h00f0: q0 = 16'h2700; // 0x01e0
	13'h00f1: q0 = 16'h4e75; // 0x01e2
	13'h00f2: q0 = 16'h4e56; // 0x01e4
	13'h00f3: q0 = 16'h0000; // 0x01e6
	13'h00f4: q0 = 16'h48e7; // 0x01e8
	13'h00f5: q0 = 16'h0f00; // 0x01ea
	13'h00f6: q0 = 16'h3e2e; // 0x01ec
	13'h00f7: q0 = 16'h0008; // 0x01ee
	13'h00f8: q0 = 16'h3c2e; // 0x01f0
	13'h00f9: q0 = 16'h000a; // 0x01f2
	13'h00fa: q0 = 16'h3a07; // 0x01f4
	13'h00fb: q0 = 16'hba46; // 0x01f6
	13'h00fc: q0 = 16'h6e20; // 0x01f8
	13'h00fd: q0 = 16'h4257; // 0x01fa
	13'h00fe: q0 = 16'h3f3c; // 0x01fc
	13'h00ff: q0 = 16'h0020; // 0x01fe
	13'h0100: q0 = 16'h3f3c; // 0x0200
	13'h0101: q0 = 16'h0064; // 0x0202
	13'h0102: q0 = 16'h3f05; // 0x0204
	13'h0103: q0 = 16'h2f3c; // 0x0206
	13'h0104: q0 = 16'h0000; // 0x0208
	13'h0105: q0 = 16'h0224; // 0x020a
	13'h0106: q0 = 16'h4eb9; // 0x020c
	13'h0107: q0 = 16'h0000; // 0x020e
	13'h0108: q0 = 16'h026c; // 0x0210
	13'h0109: q0 = 16'hdefc; // 0x0212
	13'h010a: q0 = 16'h000a; // 0x0214
	13'h010b: q0 = 16'h5245; // 0x0216
	13'h010c: q0 = 16'h60dc; // 0x0218
	13'h010d: q0 = 16'h4a9f; // 0x021a
	13'h010e: q0 = 16'h4cdf; // 0x021c
	13'h010f: q0 = 16'h00e0; // 0x021e
	13'h0110: q0 = 16'h4e5e; // 0x0220
	13'h0111: q0 = 16'h4e75; // 0x0222
	13'h0112: q0 = 16'h0000; // 0x0224
	13'h0113: q0 = 16'h4e56; // 0x0226
	13'h0114: q0 = 16'h0000; // 0x0228
	13'h0115: q0 = 16'h48e7; // 0x022a
	13'h0116: q0 = 16'h0304; // 0x022c
	13'h0117: q0 = 16'h3ebc; // 0x022e
	13'h0118: q0 = 16'h001f; // 0x0230
	13'h0119: q0 = 16'h3f3c; // 0x0232
	13'h011a: q0 = 16'h0004; // 0x0234
	13'h011b: q0 = 16'h4eb9; // 0x0236
	13'h011c: q0 = 16'h0000; // 0x0238
	13'h011d: q0 = 16'h01e4; // 0x023a
	13'h011e: q0 = 16'h4a5f; // 0x023c
	13'h011f: q0 = 16'h4247; // 0x023e
	13'h0120: q0 = 16'h2a7c; // 0x0240
	13'h0121: q0 = 16'h0001; // 0x0242
	13'h0122: q0 = 16'h8072; // 0x0244
	13'h0123: q0 = 16'hbe7c; // 0x0246
	13'h0124: q0 = 16'h0030; // 0x0248
	13'h0125: q0 = 16'h6c16; // 0x024a
	13'h0126: q0 = 16'h4255; // 0x024c
	13'h0127: q0 = 16'h426d; // 0x024e
	13'h0128: q0 = 16'h0002; // 0x0250
	13'h0129: q0 = 16'h3b7c; // 0x0252
	13'h012a: q0 = 16'h0030; // 0x0254
	13'h012b: q0 = 16'h0004; // 0x0256
	13'h012c: q0 = 16'h426d; // 0x0258
	13'h012d: q0 = 16'h0006; // 0x025a
	13'h012e: q0 = 16'h5247; // 0x025c
	13'h012f: q0 = 16'h508d; // 0x025e
	13'h0130: q0 = 16'h60e4; // 0x0260
	13'h0131: q0 = 16'h4a9f; // 0x0262
	13'h0132: q0 = 16'h4cdf; // 0x0264
	13'h0133: q0 = 16'h2080; // 0x0266
	13'h0134: q0 = 16'h4e5e; // 0x0268
	13'h0135: q0 = 16'h4e75; // 0x026a
	13'h0136: q0 = 16'h4e56; // 0x026c
	13'h0137: q0 = 16'hfffa; // 0x026e
	13'h0138: q0 = 16'h48e7; // 0x0270
	13'h0139: q0 = 16'h3f04; // 0x0272
	13'h013a: q0 = 16'h4a79; // 0x0274
	13'h013b: q0 = 16'h0001; // 0x0276
	13'h013c: q0 = 16'h7fa6; // 0x0278
	13'h013d: q0 = 16'h670c; // 0x027a
	13'h013e: q0 = 16'h302e; // 0x027c
	13'h013f: q0 = 16'h000c; // 0x027e
	13'h0140: q0 = 16'h5940; // 0x0280
	13'h0141: q0 = 16'h3d40; // 0x0282
	13'h0142: q0 = 16'h000c; // 0x0284
	13'h0143: q0 = 16'h600a; // 0x0286
	13'h0144: q0 = 16'h701f; // 0x0288
	13'h0145: q0 = 16'h906e; // 0x028a
	13'h0146: q0 = 16'h000c; // 0x028c
	13'h0147: q0 = 16'h3d40; // 0x028e
	13'h0148: q0 = 16'h000c; // 0x0290
	13'h0149: q0 = 16'h2d7c; // 0x0292
	13'h014a: q0 = 16'h0000; // 0x0294
	13'h014b: q0 = 16'h0800; // 0x0296
	13'h014c: q0 = 16'hfffa; // 0x0298
	13'h014d: q0 = 16'h202e; // 0x029a
	13'h014e: q0 = 16'hfffa; // 0x029c
	13'h014f: q0 = 16'h4281; // 0x029e
	13'h0150: q0 = 16'h720c; // 0x02a0
	13'h0151: q0 = 16'he3a0; // 0x02a2
	13'h0152: q0 = 16'h2d40; // 0x02a4
	13'h0153: q0 = 16'hfffa; // 0x02a6
	13'h0154: q0 = 16'h302e; // 0x02a8
	13'h0155: q0 = 16'h000c; // 0x02aa
	13'h0156: q0 = 16'he340; // 0x02ac
	13'h0157: q0 = 16'h48c0; // 0x02ae
	13'h0158: q0 = 16'h2a40; // 0x02b0
	13'h0159: q0 = 16'hdbee; // 0x02b2
	13'h015a: q0 = 16'hfffa; // 0x02b4
	13'h015b: q0 = 16'h2eae; // 0x02b6
	13'h015c: q0 = 16'h0008; // 0x02b8
	13'h015d: q0 = 16'h4eb9; // 0x02ba
	13'h015e: q0 = 16'h0000; // 0x02bc
	13'h015f: q0 = 16'h072e; // 0x02be
	13'h0160: q0 = 16'h3d40; // 0x02c0
	13'h0161: q0 = 16'hfffe; // 0x02c2
	13'h0162: q0 = 16'h302e; // 0x02c4
	13'h0163: q0 = 16'h0010; // 0x02c6
	13'h0164: q0 = 16'hb06e; // 0x02c8
	13'h0165: q0 = 16'hfffe; // 0x02ca
	13'h0166: q0 = 16'h6c06; // 0x02cc
	13'h0167: q0 = 16'h3d6e; // 0x02ce
	13'h0168: q0 = 16'hfffe; // 0x02d0
	13'h0169: q0 = 16'h0010; // 0x02d2
	13'h016a: q0 = 16'h0c6e; // 0x02d4
	13'h016b: q0 = 16'h0064; // 0x02d6
	13'h016c: q0 = 16'h000e; // 0x02d8
	13'h016d: q0 = 16'h6616; // 0x02da
	13'h016e: q0 = 16'h7620; // 0x02dc
	13'h016f: q0 = 16'h966e; // 0x02de
	13'h0170: q0 = 16'h0010; // 0x02e0
	13'h0171: q0 = 16'h5243; // 0x02e2
	13'h0172: q0 = 16'he243; // 0x02e4
	13'h0173: q0 = 16'h7820; // 0x02e6
	13'h0174: q0 = 16'h986e; // 0x02e8
	13'h0175: q0 = 16'hfffe; // 0x02ea
	13'h0176: q0 = 16'h5244; // 0x02ec
	13'h0177: q0 = 16'he244; // 0x02ee
	13'h0178: q0 = 16'h602c; // 0x02f0
	13'h0179: q0 = 16'h4a6e; // 0x02f2
	13'h017a: q0 = 16'h000e; // 0x02f4
	13'h017b: q0 = 16'h6c20; // 0x02f6
	13'h017c: q0 = 16'h302e; // 0x02f8
	13'h017d: q0 = 16'h000e; // 0x02fa
	13'h017e: q0 = 16'h4440; // 0x02fc
	13'h017f: q0 = 16'h3d40; // 0x02fe
	13'h0180: q0 = 16'h000e; // 0x0300
	13'h0181: q0 = 16'h362e; // 0x0302
	13'h0182: q0 = 16'h000e; // 0x0304
	13'h0183: q0 = 16'h966e; // 0x0306
	13'h0184: q0 = 16'h0010; // 0x0308
	13'h0185: q0 = 16'h5243; // 0x030a
	13'h0186: q0 = 16'h382e; // 0x030c
	13'h0187: q0 = 16'h000e; // 0x030e
	13'h0188: q0 = 16'h986e; // 0x0310
	13'h0189: q0 = 16'hfffe; // 0x0312
	13'h018a: q0 = 16'h5244; // 0x0314
	13'h018b: q0 = 16'h6006; // 0x0316
	13'h018c: q0 = 16'h362e; // 0x0318
	13'h018d: q0 = 16'h000e; // 0x031a
	13'h018e: q0 = 16'h3803; // 0x031c
	13'h018f: q0 = 16'h302e; // 0x031e
	13'h0190: q0 = 16'h0012; // 0x0320
	13'h0191: q0 = 16'hc07c; // 0x0322
	13'h0192: q0 = 16'h003f; // 0x0324
	13'h0193: q0 = 16'he140; // 0x0326
	13'h0194: q0 = 16'h3d40; // 0x0328
	13'h0195: q0 = 16'h0012; // 0x032a
	13'h0196: q0 = 16'h3e03; // 0x032c
	13'h0197: q0 = 16'h3003; // 0x032e
	13'h0198: q0 = 16'hd06e; // 0x0330
	13'h0199: q0 = 16'h0010; // 0x0332
	13'h019a: q0 = 16'hb047; // 0x0334
	13'h019b: q0 = 16'h6f64; // 0x0336
	13'h019c: q0 = 16'hbe44; // 0x0338
	13'h019d: q0 = 16'h6d0a; // 0x033a
	13'h019e: q0 = 16'h3004; // 0x033c
	13'h019f: q0 = 16'hd06e; // 0x033e
	13'h01a0: q0 = 16'hfffe; // 0x0340
	13'h01a1: q0 = 16'hb047; // 0x0342
	13'h01a2: q0 = 16'h6e04; // 0x0344
	13'h01a3: q0 = 16'h7a40; // 0x0346
	13'h01a4: q0 = 16'h6010; // 0x0348
	13'h01a5: q0 = 16'h3007; // 0x034a
	13'h01a6: q0 = 16'h9044; // 0x034c
	13'h01a7: q0 = 16'h48c0; // 0x034e
	13'h01a8: q0 = 16'hd0ae; // 0x0350
	13'h01a9: q0 = 16'h0008; // 0x0352
	13'h01aa: q0 = 16'h2040; // 0x0354
	13'h01ab: q0 = 16'h1a10; // 0x0356
	13'h01ac: q0 = 16'h4885; // 0x0358
	13'h01ad: q0 = 16'h4a79; // 0x035a
	13'h01ae: q0 = 16'h0001; // 0x035c
	13'h01af: q0 = 16'h7fa6; // 0x035e
	13'h01b0: q0 = 16'h6706; // 0x0360
	13'h01b1: q0 = 16'h7c1f; // 0x0362
	13'h01b2: q0 = 16'h9c47; // 0x0364
	13'h01b3: q0 = 16'h6002; // 0x0366
	13'h01b4: q0 = 16'h3c07; // 0x0368
	13'h01b5: q0 = 16'h4a46; // 0x036a
	13'h01b6: q0 = 16'h6606; // 0x036c
	13'h01b7: q0 = 16'h3c3c; // 0x036e
	13'h01b8: q0 = 16'h03e0; // 0x0370
	13'h01b9: q0 = 16'h6004; // 0x0372
	13'h01ba: q0 = 16'h5346; // 0x0374
	13'h01bb: q0 = 16'heb46; // 0x0376
	13'h01bc: q0 = 16'h3006; // 0x0378
	13'h01bd: q0 = 16'he340; // 0x037a
	13'h01be: q0 = 16'h48c0; // 0x037c
	13'h01bf: q0 = 16'hd08d; // 0x037e
	13'h01c0: q0 = 16'h2040; // 0x0380
	13'h01c1: q0 = 16'h3205; // 0x0382
	13'h01c2: q0 = 16'hc27c; // 0x0384
	13'h01c3: q0 = 16'h0100; // 0x0386
	13'h01c4: q0 = 16'hef41; // 0x0388
	13'h01c5: q0 = 16'h3405; // 0x038a
	13'h01c6: q0 = 16'hc47c; // 0x038c
	13'h01c7: q0 = 16'h00ff; // 0x038e
	13'h01c8: q0 = 16'h8242; // 0x0390
	13'h01c9: q0 = 16'h826e; // 0x0392
	13'h01ca: q0 = 16'h0012; // 0x0394
	13'h01cb: q0 = 16'h3081; // 0x0396
	13'h01cc: q0 = 16'h5247; // 0x0398
	13'h01cd: q0 = 16'h6092; // 0x039a
	13'h01ce: q0 = 16'h4a9f; // 0x039c
	13'h01cf: q0 = 16'h4cdf; // 0x039e
	13'h01d0: q0 = 16'h20f8; // 0x03a0
	13'h01d1: q0 = 16'h4e5e; // 0x03a2
	13'h01d2: q0 = 16'h4e75; // 0x03a4
	13'h01d3: q0 = 16'h4e56; // 0x03a6
	13'h01d4: q0 = 16'hfff6; // 0x03a8
	13'h01d5: q0 = 16'h48e7; // 0x03aa
	13'h01d6: q0 = 16'h0300; // 0x03ac
	13'h01d7: q0 = 16'h4eb9; // 0x03ae
	13'h01d8: q0 = 16'h0000; // 0x03b0
	13'h01d9: q0 = 16'h0226; // 0x03b2
	13'h01da: q0 = 16'h4279; // 0x03b4
	13'h01db: q0 = 16'h0001; // 0x03b6
	13'h01dc: q0 = 16'h7fa6; // 0x03b8
	13'h01dd: q0 = 16'h4257; // 0x03ba
	13'h01de: q0 = 16'h4267; // 0x03bc
	13'h01df: q0 = 16'h3f3c; // 0x03be
	13'h01e0: q0 = 16'h0001; // 0x03c0
	13'h01e1: q0 = 16'h3f3c; // 0x03c2
	13'h01e2: q0 = 16'h001f; // 0x03c4
	13'h01e3: q0 = 16'h2f3c; // 0x03c6
	13'h01e4: q0 = 16'h0000; // 0x03c8
	13'h01e5: q0 = 16'h0484; // 0x03ca
	13'h01e6: q0 = 16'h4eb9; // 0x03cc
	13'h01e7: q0 = 16'h0000; // 0x03ce
	13'h01e8: q0 = 16'h026c; // 0x03d0
	13'h01e9: q0 = 16'hdefc; // 0x03d2
	13'h01ea: q0 = 16'h000a; // 0x03d4
	13'h01eb: q0 = 16'h4a79; // 0x03d6
	13'h01ec: q0 = 16'h0001; // 0x03d8
	13'h01ed: q0 = 16'h7ba6; // 0x03da
	13'h01ee: q0 = 16'h6620; // 0x03dc
	13'h01ef: q0 = 16'h4257; // 0x03de
	13'h01f0: q0 = 16'h4267; // 0x03e0
	13'h01f1: q0 = 16'h3f3c; // 0x03e2
	13'h01f2: q0 = 16'h0001; // 0x03e4
	13'h01f3: q0 = 16'h3f3c; // 0x03e6
	13'h01f4: q0 = 16'h001e; // 0x03e8
	13'h01f5: q0 = 16'h2f3c; // 0x03ea
	13'h01f6: q0 = 16'h0000; // 0x03ec
	13'h01f7: q0 = 16'h048b; // 0x03ee
	13'h01f8: q0 = 16'h4eb9; // 0x03f0
	13'h01f9: q0 = 16'h0000; // 0x03f2
	13'h01fa: q0 = 16'h026c; // 0x03f4
	13'h01fb: q0 = 16'hdefc; // 0x03f6
	13'h01fc: q0 = 16'h000a; // 0x03f8
	13'h01fd: q0 = 16'h6000; // 0x03fa
	13'h01fe: q0 = 16'h007e; // 0x03fc
	13'h01ff: q0 = 16'h4247; // 0x03fe
	13'h0200: q0 = 16'hbe79; // 0x0400
	13'h0201: q0 = 16'h0001; // 0x0402
	13'h0202: q0 = 16'h7ba6; // 0x0404
	13'h0203: q0 = 16'h6c62; // 0x0406
	13'h0204: q0 = 16'h2ebc; // 0x0408
	13'h0205: q0 = 16'h0000; // 0x040a
	13'h0206: q0 = 16'h0492; // 0x040c
	13'h0207: q0 = 16'h200e; // 0x040e
	13'h0208: q0 = 16'hd0bc; // 0x0410
	13'h0209: q0 = 16'hffff; // 0x0412
	13'h020a: q0 = 16'hfff6; // 0x0414
	13'h020b: q0 = 16'h2f00; // 0x0416
	13'h020c: q0 = 16'h4eb9; // 0x0418
	13'h020d: q0 = 16'h0000; // 0x041a
	13'h020e: q0 = 16'h0750; // 0x041c
	13'h020f: q0 = 16'h4a9f; // 0x041e
	13'h0210: q0 = 16'h200e; // 0x0420
	13'h0211: q0 = 16'hd0bc; // 0x0422
	13'h0212: q0 = 16'hffff; // 0x0424
	13'h0213: q0 = 16'hfff6; // 0x0426
	13'h0214: q0 = 16'h2e80; // 0x0428
	13'h0215: q0 = 16'h3007; // 0x042a
	13'h0216: q0 = 16'he540; // 0x042c
	13'h0217: q0 = 16'h48c0; // 0x042e
	13'h0218: q0 = 16'hd0bc; // 0x0430
	13'h0219: q0 = 16'h0001; // 0x0432
	13'h021a: q0 = 16'h879e; // 0x0434
	13'h021b: q0 = 16'h2040; // 0x0436
	13'h021c: q0 = 16'h3f10; // 0x0438
	13'h021d: q0 = 16'h4eb9; // 0x043a
	13'h021e: q0 = 16'h0000; // 0x043c
	13'h021f: q0 = 16'h0798; // 0x043e
	13'h0220: q0 = 16'h4a5f; // 0x0440
	13'h0221: q0 = 16'h4257; // 0x0442
	13'h0222: q0 = 16'h4267; // 0x0444
	13'h0223: q0 = 16'h3f3c; // 0x0446
	13'h0224: q0 = 16'h0001; // 0x0448
	13'h0225: q0 = 16'h3f3c; // 0x044a
	13'h0226: q0 = 16'h001e; // 0x044c
	13'h0227: q0 = 16'h3007; // 0x044e
	13'h0228: q0 = 16'h9157; // 0x0450
	13'h0229: q0 = 16'h200e; // 0x0452
	13'h022a: q0 = 16'hd0bc; // 0x0454
	13'h022b: q0 = 16'hffff; // 0x0456
	13'h022c: q0 = 16'hfff6; // 0x0458
	13'h022d: q0 = 16'h2f00; // 0x045a
	13'h022e: q0 = 16'h4eb9; // 0x045c
	13'h022f: q0 = 16'h0000; // 0x045e
	13'h0230: q0 = 16'h026c; // 0x0460
	13'h0231: q0 = 16'hdefc; // 0x0462
	13'h0232: q0 = 16'h000a; // 0x0464
	13'h0233: q0 = 16'h5247; // 0x0466
	13'h0234: q0 = 16'h6096; // 0x0468
	13'h0235: q0 = 16'h2d79; // 0x046a
	13'h0236: q0 = 16'h0000; // 0x046c
	13'h0237: q0 = 16'h0498; // 0x046e
	13'h0238: q0 = 16'hfffc; // 0x0470
	13'h0239: q0 = 16'h206e; // 0x0472
	13'h023a: q0 = 16'hfffc; // 0x0474
	13'h023b: q0 = 16'h3e10; // 0x0476
	13'h023c: q0 = 16'h60f8; // 0x0478
	13'h023d: q0 = 16'h4a9f; // 0x047a
	13'h023e: q0 = 16'h4cdf; // 0x047c
	13'h023f: q0 = 16'h0080; // 0x047e
	13'h0240: q0 = 16'h4e5e; // 0x0480
	13'h0241: q0 = 16'h4e75; // 0x0482
	13'h0242: q0 = 16'h5241; // 0x0484
	13'h0243: q0 = 16'h4d20; // 0x0486
	13'h0244: q0 = 16'h4f4b; // 0x0488
	13'h0245: q0 = 16'h0052; // 0x048a
	13'h0246: q0 = 16'h4f4d; // 0x048c
	13'h0247: q0 = 16'h204f; // 0x048e
	13'h0248: q0 = 16'h4b00; // 0x0490
	13'h0249: q0 = 16'h524f; // 0x0492
	13'h024a: q0 = 16'h4d20; // 0x0494
	13'h024b: q0 = 16'h0000; // 0x0496
	13'h024c: q0 = 16'h0095; // 0x0498
	13'h024d: q0 = 16'h8000; // 0x049a
	13'h024e: q0 = 16'h0003; // 0x049c
	13'h024f: q0 = 16'h0080; // 0x049e
	13'h0250: q0 = 16'h0000; // 0x04a0
	13'h0251: q0 = 16'h0080; // 0x04a2
	13'h0252: q0 = 16'h07ff; // 0x04a4
	13'h0253: q0 = 16'h0001; // 0x04a6
	13'h0254: q0 = 16'h7000; // 0x04a8
	13'h0255: q0 = 16'h0001; // 0x04aa
	13'h0256: q0 = 16'h7fff; // 0x04ac
	13'h0257: q0 = 16'h0001; // 0x04ae
	13'h0258: q0 = 16'h8000; // 0x04b0
	13'h0259: q0 = 16'h0001; // 0x04b2
	13'h025a: q0 = 16'h8fff; // 0x04b4
	13'h025b: q0 = 16'h5aa5; // 0x04b6
	13'h025c: q0 = 16'h5a5a; // 0x04b8
	13'h025d: q0 = 16'ha55a; // 0x04ba
	13'h025e: q0 = 16'h5a5a; // 0x04bc
	13'h025f: q0 = 16'ha55a; // 0x04be
	13'h0260: q0 = 16'h5aa5; // 0x04c0
	13'h0261: q0 = 16'ha55a; // 0x04c2
	13'h0262: q0 = 16'ha5a5; // 0x04c4
	13'h0263: q0 = 16'h5aa5; // 0x04c6
	13'h0264: q0 = 16'h0003; // 0x04c8
	13'h0265: q0 = 16'h0000; // 0x04ca
	13'h0266: q0 = 16'h04b6; // 0x04cc
	13'h0267: q0 = 16'h0000; // 0x04ce
	13'h0268: q0 = 16'h04bc; // 0x04d0
	13'h0269: q0 = 16'h0000; // 0x04d2
	13'h026a: q0 = 16'h04c2; // 0x04d4
	13'h026b: q0 = 16'h0001; // 0x04d6
	13'h026c: q0 = 16'h4000; // 0x04d8
	13'h026d: q0 = 16'h0004; // 0x04da
	13'h026e: q0 = 16'h0000; // 0x04dc
	13'h026f: q0 = 16'h0000; // 0x04de
	13'h0270: q0 = 16'h7e0b; // 0x04e0
	13'h0271: q0 = 16'hb574; // 0x04e2
	13'h0272: q0 = 16'ha934; // 0x04e4
	13'h0273: q0 = 16'h24d8; // 0x04e6
	13'h0274: q0 = 16'h0075; // 0x04e8
	13'h0275: q0 = 16'h33fc; // 0x04ea
	13'h0276: q0 = 16'h0030; // 0x04ec
	13'h0277: q0 = 16'h0094; // 0x04ee
	13'h0278: q0 = 16'h8000; // 0x04f0
	13'h0279: q0 = 16'h323c; // 0x04f2
	13'h027a: q0 = 16'hffff; // 0x04f4
	13'h027b: q0 = 16'h4a79; // 0x04f6
	13'h027c: q0 = 16'h0095; // 0x04f8
	13'h027d: q0 = 16'h8000; // 0x04fa
`ifdef SIMULTION
 13'h0027e: 0 = 16'h4e71;
 13'h0027f: 0 = 16'h4e71;
`else
	13'h027e: q0 = 16'h51c9; // 0x04fc
	13'h027f: q0 = 16'hfff8; // 0x04fe
`endif
	13'h0280: q0 = 16'h33fc; // 0x0500
	13'h0281: q0 = 16'h0000; // 0x0502
	13'h0282: q0 = 16'h0094; // 0x0504
	13'h0283: q0 = 16'h8000; // 0x0506
	13'h0284: q0 = 16'h3639; // 0x0508
	13'h0285: q0 = 16'h0000; // 0x050a
	13'h0286: q0 = 16'h049c; // 0x050c
	13'h0287: q0 = 16'h247c; // 0x050e
	13'h0288: q0 = 16'h0000; // 0x0510
	13'h0289: q0 = 16'h049e; // 0x0512
`ifdef SIMULTION
 13'h0028a: 0 = 16'h4ef9; // 0x0514
 13'h0028b: 0 = 16'h0000; // 0x0516
 13'h0028c: 0 = 16'h0664; // 0x0518
`else
	13'h028a: q0 = 16'h6000; // 0x0514
	13'h028b: q0 = 16'h008e; // 0x0516
	13'h028c: q0 = 16'h286a; // 0x0518
`endif
	13'h028d: q0 = 16'h0004; // 0x051a
	13'h028e: q0 = 16'h3439; // 0x051c
	13'h028f: q0 = 16'h0000; // 0x051e
	13'h0290: q0 = 16'h04c8; // 0x0520
	13'h0291: q0 = 16'h227c; // 0x0522
	13'h0292: q0 = 16'h0000; // 0x0524
	13'h0293: q0 = 16'h04ca; // 0x0526
	13'h0294: q0 = 16'h6000; // 0x0528
	13'h0295: q0 = 16'h0074; // 0x052a
	13'h0296: q0 = 16'h2a51; // 0x052c
	13'h0297: q0 = 16'h2652; // 0x052e
	13'h0298: q0 = 16'h4a79; // 0x0530
	13'h0299: q0 = 16'h0095; // 0x0532
	13'h029a: q0 = 16'h8000; // 0x0534
	13'h029b: q0 = 16'h36dd; // 0x0536
	13'h029c: q0 = 16'hb7cc; // 0x0538
	13'h029d: q0 = 16'h6e10; // 0x053a
	13'h029e: q0 = 16'h36dd; // 0x053c
	13'h029f: q0 = 16'hb7cc; // 0x053e
	13'h02a0: q0 = 16'h6e0a; // 0x0540
	13'h02a1: q0 = 16'h36dd; // 0x0542
	13'h02a2: q0 = 16'hb7cc; // 0x0544
	13'h02a3: q0 = 16'h6e04; // 0x0546
	13'h02a4: q0 = 16'h5d8d; // 0x0548
	13'h02a5: q0 = 16'h60e4; // 0x054a
	13'h02a6: q0 = 16'h4a79; // 0x054c
	13'h02a7: q0 = 16'h0095; // 0x054e
	13'h02a8: q0 = 16'h8000; // 0x0550
	13'h02a9: q0 = 16'h2652; // 0x0552
	13'h02aa: q0 = 16'h2a51; // 0x0554
	13'h02ab: q0 = 16'h3815; // 0x0556
	13'h02ac: q0 = 16'h3213; // 0x0558
	13'h02ad: q0 = 16'hb841; // 0x055a
	13'h02ae: q0 = 16'h6706; // 0x055c
	13'h02af: q0 = 16'h4ef9; // 0x055e
	13'h02b0: q0 = 16'h0000; // 0x0560
	13'h02b1: q0 = 16'h05ac; // 0x0562
	13'h02b2: q0 = 16'h548d; // 0x0564
	13'h02b3: q0 = 16'h548b; // 0x0566
	13'h02b4: q0 = 16'hb7cc; // 0x0568
	13'h02b5: q0 = 16'h6e30; // 0x056a
	13'h02b6: q0 = 16'h3815; // 0x056c
	13'h02b7: q0 = 16'h3213; // 0x056e
	13'h02b8: q0 = 16'hb841; // 0x0570
	13'h02b9: q0 = 16'h6706; // 0x0572
	13'h02ba: q0 = 16'h4ef9; // 0x0574
	13'h02bb: q0 = 16'h0000; // 0x0576
	13'h02bc: q0 = 16'h05ac; // 0x0578
	13'h02bd: q0 = 16'h548d; // 0x057a
	13'h02be: q0 = 16'h548b; // 0x057c
	13'h02bf: q0 = 16'hb7cc; // 0x057e
	13'h02c0: q0 = 16'h6e1a; // 0x0580
	13'h02c1: q0 = 16'h3815; // 0x0582
	13'h02c2: q0 = 16'h3213; // 0x0584
	13'h02c3: q0 = 16'hb841; // 0x0586
	13'h02c4: q0 = 16'h6706; // 0x0588
	13'h02c5: q0 = 16'h4ef9; // 0x058a
	13'h02c6: q0 = 16'h0000; // 0x058c
	13'h02c7: q0 = 16'h05ac; // 0x058e
	13'h02c8: q0 = 16'h548d; // 0x0590
	13'h02c9: q0 = 16'h548b; // 0x0592
	13'h02ca: q0 = 16'hb7cc; // 0x0594
	13'h02cb: q0 = 16'h6e04; // 0x0596
	13'h02cc: q0 = 16'h5d8d; // 0x0598
	13'h02cd: q0 = 16'h60ba; // 0x059a
	13'h02ce: q0 = 16'h5889; // 0x059c
	13'h02cf: q0 = 16'h51ca; // 0x059e
	13'h02d0: q0 = 16'hff8c; // 0x05a0
	13'h02d1: q0 = 16'h508a; // 0x05a2
	13'h02d2: q0 = 16'h51cb; // 0x05a4
	13'h02d3: q0 = 16'hff72; // 0x05a6
	13'h02d4: q0 = 16'h6000; // 0x05a8
	13'h02d5: q0 = 16'h00ba; // 0x05aa
	13'h02d6: q0 = 16'hb344; // 0x05ac
	13'h02d7: q0 = 16'h323c; // 0x05ae
	13'h02d8: q0 = 16'h0001; // 0x05b0
	13'h02d9: q0 = 16'h3a04; // 0x05b2
	13'h02da: q0 = 16'h0245; // 0x05b4
	13'h02db: q0 = 16'h000f; // 0x05b6
	13'h02dc: q0 = 16'h6606; // 0x05b8
	13'h02dd: q0 = 16'he844; // 0x05ba
	13'h02de: q0 = 16'h5241; // 0x05bc
	13'h02df: q0 = 16'h60f2; // 0x05be
	13'h02e0: q0 = 16'hb67c; // 0x05c0
	13'h02e1: q0 = 16'h0002; // 0x05c2
	13'h02e2: q0 = 16'h664a; // 0x05c4
	13'h02e3: q0 = 16'h3801; // 0x05c6
	13'h02e4: q0 = 16'h5384; // 0x05c8
	13'h02e5: q0 = 16'h33fc; // 0x05ca
	13'h02e6: q0 = 16'h0010; // 0x05cc
	13'h02e7: q0 = 16'h0094; // 0x05ce
	13'h02e8: q0 = 16'h8000; // 0x05d0
	13'h02e9: q0 = 16'h203c; // 0x05d2
	13'h02ea: q0 = 16'h0000; // 0x05d4
	13'h02eb: q0 = 16'hffff; // 0x05d6
	13'h02ec: q0 = 16'h4a79; // 0x05d8
	13'h02ed: q0 = 16'h0095; // 0x05da
	13'h02ee: q0 = 16'h8000; // 0x05dc
`ifdef SIMULTION
	13'h02ef: q0 = 16'h4e71; // 0x05de
	13'h02f0: q0 = 16'h4e71; // 0x05e0
`else
	13'h02ef: q0 = 16'h51c8; // 0x05de
	13'h02f0: q0 = 16'hfff8; // 0x05e0
`endif
	13'h02f1: q0 = 16'h33fc; // 0x05e2
	13'h02f2: q0 = 16'h0000; // 0x05e4
	13'h02f3: q0 = 16'h0094; // 0x05e6
	13'h02f4: q0 = 16'h8000; // 0x05e8
	13'h02f5: q0 = 16'h203c; // 0x05ea
	13'h02f6: q0 = 16'h0000; // 0x05ec
	13'h02f7: q0 = 16'hffff; // 0x05ee
	13'h02f8: q0 = 16'h4a79; // 0x05f0
	13'h02f9: q0 = 16'h0095; // 0x05f2
	13'h02fa: q0 = 16'h8000; // 0x05f4
`ifdef SIMULTION
	13'h02fb: q0 = 16'h4e71; // 0x05f6
	13'h02fc: q0 = 16'h4e71; // 0x05f8
`else
	13'h02fb: q0 = 16'h51c8; // 0x05f6
	13'h02fc: q0 = 16'hfff8; // 0x05f8
`endif
	13'h02fd: q0 = 16'h51cc; // 0x05fa
	13'h02fe: q0 = 16'hffce; // 0x05fc
	13'h02ff: q0 = 16'h203c; // 0x05fe
	13'h0300: q0 = 16'h0001; // 0x0600
	13'h0301: q0 = 16'hffff; // 0x0602
	13'h0302: q0 = 16'h4a79; // 0x0604
	13'h0303: q0 = 16'h0095; // 0x0606
	13'h0304: q0 = 16'h8000; // 0x0608
`ifdef SIMULTION
	13'h0305: q0 = 16'h4e71; // 0x060a
	13'h0306: q0 = 16'h4e71; // 0x060c
`else
	13'h0305: q0 = 16'h51c8; // 0x060a
	13'h0306: q0 = 16'hfff8; // 0x060c
`endif
	13'h0307: q0 = 16'h60b6; // 0x060e
	13'h0308: q0 = 16'h33fc; // 0x0610
	13'h0309: q0 = 16'h0010; // 0x0612
	13'h030a: q0 = 16'h0094; // 0x0614
	13'h030b: q0 = 16'h8000; // 0x0616
	13'h030c: q0 = 16'hb27c; // 0x0618
	13'h030d: q0 = 16'h0003; // 0x061a
	13'h030e: q0 = 16'h6d02; // 0x061c
	13'h030f: q0 = 16'h5443; // 0x061e
	13'h0310: q0 = 16'h383c; // 0x0620
	13'h0311: q0 = 16'h03ff; // 0x0622
	13'h0312: q0 = 16'h227c; // 0x0624
	13'h0313: q0 = 16'h0080; // 0x0626
	13'h0314: q0 = 16'h0000; // 0x0628
	13'h0315: q0 = 16'h32fc; // 0x062a
	13'h0316: q0 = 16'h0020; // 0x062c
	13'h0317: q0 = 16'h51cc; // 0x062e
	13'h0318: q0 = 16'hfffa; // 0x0630
	13'h0319: q0 = 16'h227c; // 0x0632
	13'h031a: q0 = 16'h0080; // 0x0634
	13'h031b: q0 = 16'h0000; // 0x0636
	13'h031c: q0 = 16'h32bc; // 0x0638
	13'h031d: q0 = 16'h0052; // 0x063a
	13'h031e: q0 = 16'hd3fc; // 0x063c
	13'h031f: q0 = 16'h0000; // 0x063e
	13'h0320: q0 = 16'h0040; // 0x0640
	13'h0321: q0 = 16'h32bc; // 0x0642
	13'h0322: q0 = 16'h0041; // 0x0644
	13'h0323: q0 = 16'hd3fc; // 0x0646
	13'h0324: q0 = 16'h0000; // 0x0648
	13'h0325: q0 = 16'h0040; // 0x064a
	13'h0326: q0 = 16'h32bc; // 0x064c
	13'h0327: q0 = 16'h004d; // 0x064e
	13'h0328: q0 = 16'hd3fc; // 0x0650
	13'h0329: q0 = 16'h0000; // 0x0652
	13'h032a: q0 = 16'h0080; // 0x0654
	13'h032b: q0 = 16'hd67c; // 0x0656
	13'h032c: q0 = 16'h0030; // 0x0658
	13'h032d: q0 = 16'h3283; // 0x065a
	13'h032e: q0 = 16'h4a79; // 0x065c
	13'h032f: q0 = 16'h0095; // 0x065e
	13'h0330: q0 = 16'h8000; // 0x0660
	13'h0331: q0 = 16'h60f8; // 0x0662
	13'h0332: q0 = 16'h4e71; // 0x0664
	13'h0333: q0 = 16'h33fc; // 0x0666
	13'h0334: q0 = 16'h0020; // 0x0668
	13'h0335: q0 = 16'h0001; // 0x066a
	13'h0336: q0 = 16'h861e; // 0x066c
	13'h0337: q0 = 16'h33f9; // 0x066e
	13'h0338: q0 = 16'h0001; // 0x0670
	13'h0339: q0 = 16'h861e; // 0x0672
	13'h033a: q0 = 16'h0094; // 0x0674
	13'h033b: q0 = 16'h8000; // 0x0676
	13'h033c: q0 = 16'h207c; // 0x0678
	13'h033d: q0 = 16'h0001; // 0x067a
	13'h033e: q0 = 16'h879c; // 0x067c
	13'h033f: q0 = 16'h4280; // 0x067e
	13'h0340: q0 = 16'h227c; // 0x0680
	13'h0341: q0 = 16'h0000; // 0x0682
	13'h0342: q0 = 16'h04e0; // 0x0684
	13'h0343: q0 = 16'h4281; // 0x0686
`ifdef SIMULTION
 13'h00344: 0 = 16'h4241; // 0x0688
 13'h00345: 0 = 16'h4e71; // 0x068a
 13'h00346: 0 = 16'h4e71; // 0x068c
`else
	13'h0344: q0 = 16'hb279; // 0x0688
	13'h0345: q0 = 16'h0000; // 0x068a
	13'h0346: q0 = 16'h04d6; // 0x068c
`endif
	13'h0347: q0 = 16'h6c00; // 0x068e
	13'h0348: q0 = 16'h0076; // 0x0690
	13'h0349: q0 = 16'h2a01; // 0x0692
	13'h034a: q0 = 16'he345; // 0x0694
	13'h034b: q0 = 16'he345; // 0x0696
	13'h034c: q0 = 16'h2a7c; // 0x0698
	13'h034d: q0 = 16'h0000; // 0x069a
	13'h034e: q0 = 16'h04dc; // 0x069c
	13'h034f: q0 = 16'hdbc5; // 0x069e
	13'h0350: q0 = 16'h2455; // 0x06a0
	13'h0351: q0 = 16'he245; // 0x06a2
	13'h0352: q0 = 16'h4242; // 0x06a4
	13'h0353: q0 = 16'h4a79; // 0x06a6
	13'h0354: q0 = 16'h0095; // 0x06a8
	13'h0355: q0 = 16'h8000; // 0x06aa
	13'h0356: q0 = 16'h2a7c; // 0x06ac
	13'h0357: q0 = 16'h0000; // 0x06ae
	13'h0358: q0 = 16'h04da; // 0x06b0
	13'h0359: q0 = 16'hdbc5; // 0x06b2
	13'h035a: q0 = 16'hb455; // 0x06b4
	13'h035b: q0 = 16'h6c4a; // 0x06b6
	13'h035c: q0 = 16'h4203; // 0x06b8
	13'h035d: q0 = 16'h4204; // 0x06ba
	13'h035e: q0 = 16'h264a; // 0x06bc
	13'h035f: q0 = 16'h2a7c; // 0x06be
	13'h0360: q0 = 16'h0000; // 0x06c0
	13'h0361: q0 = 16'h04d8; // 0x06c2
	13'h0362: q0 = 16'hdbc5; // 0x06c4
	13'h0363: q0 = 16'h3c15; // 0x06c6
	13'h0364: q0 = 16'h48c6; // 0x06c8
	13'h0365: q0 = 16'hd7c6; // 0x06ca
	13'h0366: q0 = 16'h4246; // 0x06cc
	13'h0367: q0 = 16'hb5cb; // 0x06ce
	13'h0368: q0 = 16'h6c06; // 0x06d0
	13'h0369: q0 = 16'hd61a; // 0x06d2
	13'h036a: q0 = 16'hd81a; // 0x06d4
	13'h036b: q0 = 16'h60f6; // 0x06d6
	13'h036c: q0 = 16'hb619; // 0x06d8
	13'h036d: q0 = 16'h670e; // 0x06da
	13'h036e: q0 = 16'h0c40; // 0x06dc
	13'h036f: q0 = 16'h0010; // 0x06de
	13'h0370: q0 = 16'h6c08; // 0x06e0
	13'h0371: q0 = 16'h30c1; // 0x06e2
	13'h0372: q0 = 16'h3082; // 0x06e4
	13'h0373: q0 = 16'he1d8; // 0x06e6
	13'h0374: q0 = 16'h5240; // 0x06e8
	13'h0375: q0 = 16'hb819; // 0x06ea
	13'h0376: q0 = 16'h6710; // 0x06ec
	13'h0377: q0 = 16'h0c40; // 0x06ee
	13'h0378: q0 = 16'h0010; // 0x06f0
	13'h0379: q0 = 16'h6c0a; // 0x06f2
	13'h037a: q0 = 16'h30c1; // 0x06f4
	13'h037b: q0 = 16'h3082; // 0x06f6
	13'h037c: q0 = 16'he1d0; // 0x06f8
	13'h037d: q0 = 16'h5258; // 0x06fa
	13'h037e: q0 = 16'h5240; // 0x06fc
	13'h037f: q0 = 16'h5242; // 0x06fe
	13'h0380: q0 = 16'h60a4; // 0x0700
	13'h0381: q0 = 16'h5241; // 0x0702
	13'h0382: q0 = 16'h6082; // 0x0704
`ifdef SIMULTION
 13'h00383: 0 = 16'h4240; // 0x0706
`else
	13'h0383: q0 = 16'h4a40; // 0x0706
`endif
	13'h0384: q0 = 16'h6612; // 0x0708
	13'h0385: q0 = 16'h0279; // 0x070a
	13'h0386: q0 = 16'hffdf; // 0x070c
	13'h0387: q0 = 16'h0001; // 0x070e
	13'h0388: q0 = 16'h861e; // 0x0710
	13'h0389: q0 = 16'h33f9; // 0x0712
	13'h038a: q0 = 16'h0001; // 0x0714
	13'h038b: q0 = 16'h861e; // 0x0716
	13'h038c: q0 = 16'h0094; // 0x0718
	13'h038d: q0 = 16'h8000; // 0x071a
	13'h038e: q0 = 16'h33c0; // 0x071c
	13'h038f: q0 = 16'h0001; // 0x071e
	13'h0390: q0 = 16'h7ba6; // 0x0720
	13'h0391: q0 = 16'h4eb9; // 0x0722
	13'h0392: q0 = 16'h0000; // 0x0724
	13'h0393: q0 = 16'h03a6; // 0x0726
	13'h0394: q0 = 16'h4ef9; // 0x0728
	13'h0395: q0 = 16'h0000; // 0x072a
	13'h0396: q0 = 16'h00d4; // 0x072c
	13'h0397: q0 = 16'h4e56; // 0x072e
	13'h0398: q0 = 16'h0000; // 0x0730
	13'h0399: q0 = 16'h48e7; // 0x0732
	13'h039a: q0 = 16'h0304; // 0x0734
	13'h039b: q0 = 16'h2a6e; // 0x0736
	13'h039c: q0 = 16'h0008; // 0x0738
	13'h039d: q0 = 16'h4247; // 0x073a
	13'h039e: q0 = 16'h4a1d; // 0x073c
	13'h039f: q0 = 16'h6704; // 0x073e
	13'h03a0: q0 = 16'h5247; // 0x0740
	13'h03a1: q0 = 16'h60f8; // 0x0742
	13'h03a2: q0 = 16'h3007; // 0x0744
	13'h03a3: q0 = 16'h4a9f; // 0x0746
	13'h03a4: q0 = 16'h4cdf; // 0x0748
	13'h03a5: q0 = 16'h2080; // 0x074a
	13'h03a6: q0 = 16'h4e5e; // 0x074c
	13'h03a7: q0 = 16'h4e75; // 0x074e
	13'h03a8: q0 = 16'h4e56; // 0x0750
	13'h03a9: q0 = 16'h0000; // 0x0752
	13'h03aa: q0 = 16'h48e7; // 0x0754
	13'h03ab: q0 = 16'h010c; // 0x0756
	13'h03ac: q0 = 16'h2a6e; // 0x0758
	13'h03ad: q0 = 16'h0008; // 0x075a
	13'h03ae: q0 = 16'h286e; // 0x075c
	13'h03af: q0 = 16'h000c; // 0x075e
	13'h03b0: q0 = 16'h1adc; // 0x0760
	13'h03b1: q0 = 16'h6702; // 0x0762
	13'h03b2: q0 = 16'h60fa; // 0x0764
	13'h03b3: q0 = 16'h4a9f; // 0x0766
	13'h03b4: q0 = 16'h4cdf; // 0x0768
	13'h03b5: q0 = 16'h3000; // 0x076a
	13'h03b6: q0 = 16'h4e5e; // 0x076c
	13'h03b7: q0 = 16'h4e75; // 0x076e
	13'h03b8: q0 = 16'h4e56; // 0x0770
	13'h03b9: q0 = 16'h0000; // 0x0772
	13'h03ba: q0 = 16'h48e7; // 0x0774
	13'h03bb: q0 = 16'h010c; // 0x0776
	13'h03bc: q0 = 16'h2a6e; // 0x0778
	13'h03bd: q0 = 16'h0008; // 0x077a
	13'h03be: q0 = 16'h286e; // 0x077c
	13'h03bf: q0 = 16'h000c; // 0x077e
	13'h03c0: q0 = 16'h4a15; // 0x0780
	13'h03c1: q0 = 16'h6704; // 0x0782
	13'h03c2: q0 = 16'h528d; // 0x0784
	13'h03c3: q0 = 16'h60f8; // 0x0786
	13'h03c4: q0 = 16'h1adc; // 0x0788
	13'h03c5: q0 = 16'h6702; // 0x078a
	13'h03c6: q0 = 16'h60fa; // 0x078c
	13'h03c7: q0 = 16'h4a9f; // 0x078e
	13'h03c8: q0 = 16'h4cdf; // 0x0790
	13'h03c9: q0 = 16'h3000; // 0x0792
	13'h03ca: q0 = 16'h4e5e; // 0x0794
	13'h03cb: q0 = 16'h4e75; // 0x0796
	13'h03cc: q0 = 16'h4e56; // 0x0798
	13'h03cd: q0 = 16'hfffc; // 0x079a
	13'h03ce: q0 = 16'h48e7; // 0x079c
	13'h03cf: q0 = 16'h0104; // 0x079e
	13'h03d0: q0 = 16'h2a6e; // 0x07a0
	13'h03d1: q0 = 16'h000a; // 0x07a2
	13'h03d2: q0 = 16'h4a15; // 0x07a4
	13'h03d3: q0 = 16'h6704; // 0x07a6
	13'h03d4: q0 = 16'h528d; // 0x07a8
	13'h03d5: q0 = 16'h60f8; // 0x07aa
	13'h03d6: q0 = 16'h2d4d; // 0x07ac
	13'h03d7: q0 = 16'hfffc; // 0x07ae
	13'h03d8: q0 = 16'h2eae; // 0x07b0
	13'h03d9: q0 = 16'hfffc; // 0x07b2
	13'h03da: q0 = 16'h3f2e; // 0x07b4
	13'h03db: q0 = 16'h0008; // 0x07b6
	13'h03dc: q0 = 16'h616e; // 0x07b8
	13'h03dd: q0 = 16'h4a5f; // 0x07ba
	13'h03de: q0 = 16'h4a9f; // 0x07bc
	13'h03df: q0 = 16'h4cdf; // 0x07be
	13'h03e0: q0 = 16'h2000; // 0x07c0
	13'h03e1: q0 = 16'h4e5e; // 0x07c2
	13'h03e2: q0 = 16'h4e75; // 0x07c4
	13'h03e3: q0 = 16'h4e56; // 0x07c6
	13'h03e4: q0 = 16'hfffc; // 0x07c8
	13'h03e5: q0 = 16'h48e7; // 0x07ca
	13'h03e6: q0 = 16'h0104; // 0x07cc
	13'h03e7: q0 = 16'h2a6e; // 0x07ce
	13'h03e8: q0 = 16'h000c; // 0x07d0
	13'h03e9: q0 = 16'h4a15; // 0x07d2
	13'h03ea: q0 = 16'h6704; // 0x07d4
	13'h03eb: q0 = 16'h528d; // 0x07d6
	13'h03ec: q0 = 16'h60f8; // 0x07d8
	13'h03ed: q0 = 16'h2d4d; // 0x07da
	13'h03ee: q0 = 16'hfffc; // 0x07dc
	13'h03ef: q0 = 16'h2eae; // 0x07de
	13'h03f0: q0 = 16'hfffc; // 0x07e0
	13'h03f1: q0 = 16'h2f2e; // 0x07e2
	13'h03f2: q0 = 16'h0008; // 0x07e4
	13'h03f3: q0 = 16'h6100; // 0x07e6
	13'h03f4: q0 = 16'h00aa; // 0x07e8
	13'h03f5: q0 = 16'h4a9f; // 0x07ea
	13'h03f6: q0 = 16'h4a9f; // 0x07ec
	13'h03f7: q0 = 16'h4cdf; // 0x07ee
	13'h03f8: q0 = 16'h2000; // 0x07f0
	13'h03f9: q0 = 16'h4e5e; // 0x07f2
	13'h03fa: q0 = 16'h4e75; // 0x07f4
	13'h03fb: q0 = 16'h4e56; // 0x07f6
	13'h03fc: q0 = 16'h0000; // 0x07f8
	13'h03fd: q0 = 16'h48e7; // 0x07fa
	13'h03fe: q0 = 16'h030c; // 0x07fc
	13'h03ff: q0 = 16'h2a6e; // 0x07fe
	13'h0400: q0 = 16'h0008; // 0x0800
	13'h0401: q0 = 16'h284d; // 0x0802
	13'h0402: q0 = 16'h4a14; // 0x0804
	13'h0403: q0 = 16'h6704; // 0x0806
	13'h0404: q0 = 16'h528c; // 0x0808
	13'h0405: q0 = 16'h60f8; // 0x080a
	13'h0406: q0 = 16'h538c; // 0x080c
	13'h0407: q0 = 16'hbbcc; // 0x080e
	13'h0408: q0 = 16'h640c; // 0x0810
	13'h0409: q0 = 16'h1e15; // 0x0812
	13'h040a: q0 = 16'h1a94; // 0x0814
	13'h040b: q0 = 16'h1887; // 0x0816
	13'h040c: q0 = 16'h528d; // 0x0818
	13'h040d: q0 = 16'h538c; // 0x081a
	13'h040e: q0 = 16'h60f0; // 0x081c
	13'h040f: q0 = 16'h4a9f; // 0x081e
	13'h0410: q0 = 16'h4cdf; // 0x0820
	13'h0411: q0 = 16'h3080; // 0x0822
	13'h0412: q0 = 16'h4e5e; // 0x0824
	13'h0413: q0 = 16'h4e75; // 0x0826
	13'h0414: q0 = 16'h4e56; // 0x0828
	13'h0415: q0 = 16'hfffa; // 0x082a
	13'h0416: q0 = 16'h48e7; // 0x082c
	13'h0417: q0 = 16'h0304; // 0x082e
	13'h0418: q0 = 16'h3e2e; // 0x0830
	13'h0419: q0 = 16'h0008; // 0x0832
	13'h041a: q0 = 16'h2a6e; // 0x0834
	13'h041b: q0 = 16'h000a; // 0x0836
	13'h041c: q0 = 16'h2d4d; // 0x0838
	13'h041d: q0 = 16'hfffa; // 0x083a
	13'h041e: q0 = 16'h3d47; // 0x083c
	13'h041f: q0 = 16'hfffe; // 0x083e
	13'h0420: q0 = 16'h6c06; // 0x0840
	13'h0421: q0 = 16'h3007; // 0x0842
	13'h0422: q0 = 16'h4440; // 0x0844
	13'h0423: q0 = 16'h3e00; // 0x0846
	13'h0424: q0 = 16'hbe7c; // 0x0848
	13'h0425: q0 = 16'h000a; // 0x084a
	13'h0426: q0 = 16'h6c0a; // 0x084c
	13'h0427: q0 = 16'h3007; // 0x084e
	13'h0428: q0 = 16'hd07c; // 0x0850
	13'h0429: q0 = 16'h0030; // 0x0852
	13'h042a: q0 = 16'h1ac0; // 0x0854
	13'h042b: q0 = 16'h601c; // 0x0856
	13'h042c: q0 = 16'h3007; // 0x0858
	13'h042d: q0 = 16'h48c0; // 0x085a
	13'h042e: q0 = 16'h81fc; // 0x085c
	13'h042f: q0 = 16'h000a; // 0x085e
	13'h0430: q0 = 16'h4840; // 0x0860
	13'h0431: q0 = 16'hd07c; // 0x0862
	13'h0432: q0 = 16'h0030; // 0x0864
	13'h0433: q0 = 16'h1ac0; // 0x0866
	13'h0434: q0 = 16'h3007; // 0x0868
	13'h0435: q0 = 16'h48c0; // 0x086a
	13'h0436: q0 = 16'h81fc; // 0x086c
	13'h0437: q0 = 16'h000a; // 0x086e
	13'h0438: q0 = 16'h3e00; // 0x0870
	13'h0439: q0 = 16'h6ee4; // 0x0872
	13'h043a: q0 = 16'h4a6e; // 0x0874
	13'h043b: q0 = 16'hfffe; // 0x0876
	13'h043c: q0 = 16'h6c04; // 0x0878
	13'h043d: q0 = 16'h1afc; // 0x087a
	13'h043e: q0 = 16'h002d; // 0x087c
	13'h043f: q0 = 16'h4215; // 0x087e
	13'h0440: q0 = 16'h2eae; // 0x0880
	13'h0441: q0 = 16'hfffa; // 0x0882
	13'h0442: q0 = 16'h6100; // 0x0884
	13'h0443: q0 = 16'hff70; // 0x0886
	13'h0444: q0 = 16'h4a9f; // 0x0888
	13'h0445: q0 = 16'h4cdf; // 0x088a
	13'h0446: q0 = 16'h2080; // 0x088c
	13'h0447: q0 = 16'h4e5e; // 0x088e
	13'h0448: q0 = 16'h4e75; // 0x0890
	13'h0449: q0 = 16'h4e56; // 0x0892
	13'h044a: q0 = 16'hfff8; // 0x0894
	13'h044b: q0 = 16'h48e7; // 0x0896
	13'h044c: q0 = 16'h0704; // 0x0898
	13'h044d: q0 = 16'h2e2e; // 0x089a
	13'h044e: q0 = 16'h0008; // 0x089c
	13'h044f: q0 = 16'h2a6e; // 0x089e
	13'h0450: q0 = 16'h000c; // 0x08a0
	13'h0451: q0 = 16'h2d4d; // 0x08a2
	13'h0452: q0 = 16'hfff8; // 0x08a4
	13'h0453: q0 = 16'h2d47; // 0x08a6
	13'h0454: q0 = 16'hfffc; // 0x08a8
	13'h0455: q0 = 16'h6c06; // 0x08aa
	13'h0456: q0 = 16'h2007; // 0x08ac
	13'h0457: q0 = 16'h4480; // 0x08ae
	13'h0458: q0 = 16'h2e00; // 0x08b0
	13'h0459: q0 = 16'h2f39; // 0x08b2
	13'h045a: q0 = 16'h0000; // 0x08b4
	13'h045b: q0 = 16'hc100; // 0x08b6
	13'h045c: q0 = 16'h2f07; // 0x08b8
	13'h045d: q0 = 16'h4eb9; // 0x08ba
	13'h045e: q0 = 16'h0000; // 0x08bc
	13'h045f: q0 = 16'h79ac; // 0x08be
	13'h0460: q0 = 16'hbf8f; // 0x08c0
	13'h0461: q0 = 16'h2c00; // 0x08c2
	13'h0462: q0 = 16'h2f39; // 0x08c4
	13'h0463: q0 = 16'h0000; // 0x08c6
	13'h0464: q0 = 16'hc100; // 0x08c8
	13'h0465: q0 = 16'h2f06; // 0x08ca
	13'h0466: q0 = 16'h4eb9; // 0x08cc
	13'h0467: q0 = 16'h0000; // 0x08ce
	13'h0468: q0 = 16'h7a50; // 0x08d0
	13'h0469: q0 = 16'hbf8f; // 0x08d2
	13'h046a: q0 = 16'h2f00; // 0x08d4
	13'h046b: q0 = 16'h2007; // 0x08d6
	13'h046c: q0 = 16'h221f; // 0x08d8
	13'h046d: q0 = 16'h9081; // 0x08da
	13'h046e: q0 = 16'hd0bc; // 0x08dc
	13'h046f: q0 = 16'h0000; // 0x08de
	13'h0470: q0 = 16'h0030; // 0x08e0
	13'h0471: q0 = 16'h1ac0; // 0x08e2
	13'h0472: q0 = 16'h2e06; // 0x08e4
	13'h0473: q0 = 16'h4a87; // 0x08e6
	13'h0474: q0 = 16'h6ec8; // 0x08e8
	13'h0475: q0 = 16'h4aae; // 0x08ea
	13'h0476: q0 = 16'hfffc; // 0x08ec
	13'h0477: q0 = 16'h6c04; // 0x08ee
	13'h0478: q0 = 16'h1afc; // 0x08f0
	13'h0479: q0 = 16'h002d; // 0x08f2
	13'h047a: q0 = 16'h4215; // 0x08f4
	13'h047b: q0 = 16'h2eae; // 0x08f6
	13'h047c: q0 = 16'hfff8; // 0x08f8
	13'h047d: q0 = 16'h6100; // 0x08fa
	13'h047e: q0 = 16'hfefa; // 0x08fc
	13'h047f: q0 = 16'h4a9f; // 0x08fe
	13'h0480: q0 = 16'h4cdf; // 0x0900
	13'h0481: q0 = 16'h20c0; // 0x0902
	13'h0482: q0 = 16'h4e5e; // 0x0904
	13'h0483: q0 = 16'h4e75; // 0x0906
	13'h0484: q0 = 16'h4e56; // 0x0908
	13'h0485: q0 = 16'h0000; // 0x090a
	13'h0486: q0 = 16'h48e7; // 0x090c
	13'h0487: q0 = 16'h0304; // 0x090e
	13'h0488: q0 = 16'h4247; // 0x0910
	13'h0489: q0 = 16'h2eae; // 0x0912
	13'h048a: q0 = 16'h000c; // 0x0914
	13'h048b: q0 = 16'h6100; // 0x0916
	13'h048c: q0 = 16'hfede; // 0x0918
	13'h048d: q0 = 16'h2eae; // 0x091a
	13'h048e: q0 = 16'h0008; // 0x091c
	13'h048f: q0 = 16'h6100; // 0x091e
	13'h0490: q0 = 16'hfed6; // 0x0920
	13'h0491: q0 = 16'h2a6e; // 0x0922
	13'h0492: q0 = 16'h0008; // 0x0924
	13'h0493: q0 = 16'h4a15; // 0x0926
	13'h0494: q0 = 16'h660e; // 0x0928
	13'h0495: q0 = 16'h202e; // 0x092a
	13'h0496: q0 = 16'h000c; // 0x092c
	13'h0497: q0 = 16'h2040; // 0x092e
	13'h0498: q0 = 16'h4a10; // 0x0930
	13'h0499: q0 = 16'h6604; // 0x0932
	13'h049a: q0 = 16'h4a47; // 0x0934
	13'h049b: q0 = 16'h6758; // 0x0936
	13'h049c: q0 = 16'h4a15; // 0x0938
	13'h049d: q0 = 16'h660e; // 0x093a
	13'h049e: q0 = 16'h2ebc; // 0x093c
	13'h049f: q0 = 16'h0000; // 0x093e
	13'h04a0: q0 = 16'hc104; // 0x0940
	13'h04a1: q0 = 16'h2f0d; // 0x0942
	13'h04a2: q0 = 16'h6100; // 0x0944
	13'h04a3: q0 = 16'hfe2a; // 0x0946
	13'h04a4: q0 = 16'h4a9f; // 0x0948
	13'h04a5: q0 = 16'h202e; // 0x094a
	13'h04a6: q0 = 16'h000c; // 0x094c
	13'h04a7: q0 = 16'h2040; // 0x094e
	13'h04a8: q0 = 16'h4a10; // 0x0950
	13'h04a9: q0 = 16'h6714; // 0x0952
	13'h04aa: q0 = 16'h202e; // 0x0954
	13'h04ab: q0 = 16'h000c; // 0x0956
	13'h04ac: q0 = 16'h2040; // 0x0958
	13'h04ad: q0 = 16'h1010; // 0x095a
	13'h04ae: q0 = 16'h4880; // 0x095c
	13'h04af: q0 = 16'hd07c; // 0x095e
	13'h04b0: q0 = 16'hffd0; // 0x0960
	13'h04b1: q0 = 16'h1215; // 0x0962
	13'h04b2: q0 = 16'hd200; // 0x0964
	13'h04b3: q0 = 16'h1a81; // 0x0966
	13'h04b4: q0 = 16'h4a47; // 0x0968
	13'h04b5: q0 = 16'h6702; // 0x096a
	13'h04b6: q0 = 16'h5215; // 0x096c
	13'h04b7: q0 = 16'h0c15; // 0x096e
	13'h04b8: q0 = 16'h0039; // 0x0970
	13'h04b9: q0 = 16'h6f08; // 0x0972
	13'h04ba: q0 = 16'h0415; // 0x0974
	13'h04bb: q0 = 16'h000a; // 0x0976
	13'h04bc: q0 = 16'h7e01; // 0x0978
	13'h04bd: q0 = 16'h6002; // 0x097a
	13'h04be: q0 = 16'h4247; // 0x097c
	13'h04bf: q0 = 16'h202e; // 0x097e
	13'h04c0: q0 = 16'h000c; // 0x0980
	13'h04c1: q0 = 16'h2040; // 0x0982
	13'h04c2: q0 = 16'h4a10; // 0x0984
	13'h04c3: q0 = 16'h6704; // 0x0986
	13'h04c4: q0 = 16'h52ae; // 0x0988
	13'h04c5: q0 = 16'h000c; // 0x098a
	13'h04c6: q0 = 16'h528d; // 0x098c
	13'h04c7: q0 = 16'h6096; // 0x098e
	13'h04c8: q0 = 16'h2eae; // 0x0990
	13'h04c9: q0 = 16'h0008; // 0x0992
	13'h04ca: q0 = 16'h6100; // 0x0994
	13'h04cb: q0 = 16'hfe60; // 0x0996
	13'h04cc: q0 = 16'h4a9f; // 0x0998
	13'h04cd: q0 = 16'h4cdf; // 0x099a
	13'h04ce: q0 = 16'h2080; // 0x099c
	13'h04cf: q0 = 16'h4e5e; // 0x099e
	13'h04d0: q0 = 16'h4e75; // 0x09a0
	13'h04d1: q0 = 16'h4e56; // 0x09a2
	13'h04d2: q0 = 16'hfffc; // 0x09a4
	13'h04d3: q0 = 16'h4a6e; // 0x09a6
	13'h04d4: q0 = 16'h0008; // 0x09a8
	13'h04d5: q0 = 16'h6c08; // 0x09aa
	13'h04d6: q0 = 16'h302e; // 0x09ac
	13'h04d7: q0 = 16'h0008; // 0x09ae
	13'h04d8: q0 = 16'h4440; // 0x09b0
	13'h04d9: q0 = 16'h6004; // 0x09b2
	13'h04da: q0 = 16'h302e; // 0x09b4
	13'h04db: q0 = 16'h0008; // 0x09b6
	13'h04dc: q0 = 16'h4e5e; // 0x09b8
	13'h04dd: q0 = 16'h4e75; // 0x09ba
	13'h04de: q0 = 16'h4e56; // 0x09bc
	13'h04df: q0 = 16'h0000; // 0x09be
	13'h04e0: q0 = 16'h48e7; // 0x09c0
	13'h04e1: q0 = 16'h0f0c; // 0x09c2
	13'h04e2: q0 = 16'h3e2e; // 0x09c4
	13'h04e3: q0 = 16'h0008; // 0x09c6
	13'h04e4: q0 = 16'h2a6e; // 0x09c8
	13'h04e5: q0 = 16'h000a; // 0x09ca
	13'h04e6: q0 = 16'h286e; // 0x09cc
	13'h04e7: q0 = 16'h000e; // 0x09ce
	13'h04e8: q0 = 16'h4245; // 0x09d0
	13'h04e9: q0 = 16'h4246; // 0x09d2
	13'h04ea: q0 = 16'h4a55; // 0x09d4
	13'h04eb: q0 = 16'h6c08; // 0x09d6
	13'h04ec: q0 = 16'h7a01; // 0x09d8
	13'h04ed: q0 = 16'h3015; // 0x09da
	13'h04ee: q0 = 16'h4440; // 0x09dc
	13'h04ef: q0 = 16'h3a80; // 0x09de
	13'h04f0: q0 = 16'h4a54; // 0x09e0
	13'h04f1: q0 = 16'h6c08; // 0x09e2
	13'h04f2: q0 = 16'h7c01; // 0x09e4
	13'h04f3: q0 = 16'h3014; // 0x09e6
	13'h04f4: q0 = 16'h4440; // 0x09e8
	13'h04f5: q0 = 16'h3880; // 0x09ea
	13'h04f6: q0 = 16'h3015; // 0x09ec
	13'h04f7: q0 = 16'hb047; // 0x09ee
	13'h04f8: q0 = 16'h6e06; // 0x09f0
	13'h04f9: q0 = 16'h3014; // 0x09f2
	13'h04fa: q0 = 16'hb047; // 0x09f4
	13'h04fb: q0 = 16'h6f06; // 0x09f6
	13'h04fc: q0 = 16'he0d5; // 0x09f8
	13'h04fd: q0 = 16'he0d4; // 0x09fa
	13'h04fe: q0 = 16'h60ee; // 0x09fc
	13'h04ff: q0 = 16'h4a45; // 0x09fe
	13'h0500: q0 = 16'h6706; // 0x0a00
	13'h0501: q0 = 16'h3015; // 0x0a02
	13'h0502: q0 = 16'h4440; // 0x0a04
	13'h0503: q0 = 16'h3a80; // 0x0a06
	13'h0504: q0 = 16'h4a46; // 0x0a08
	13'h0505: q0 = 16'h6706; // 0x0a0a
	13'h0506: q0 = 16'h3014; // 0x0a0c
	13'h0507: q0 = 16'h4440; // 0x0a0e
	13'h0508: q0 = 16'h3880; // 0x0a10
	13'h0509: q0 = 16'h4a9f; // 0x0a12
	13'h050a: q0 = 16'h4cdf; // 0x0a14
	13'h050b: q0 = 16'h30e0; // 0x0a16
	13'h050c: q0 = 16'h4e5e; // 0x0a18
	13'h050d: q0 = 16'h4e75; // 0x0a1a
	13'h050e: q0 = 16'h4e56; // 0x0a1c
	13'h050f: q0 = 16'h0000; // 0x0a1e
	13'h0510: q0 = 16'h48e7; // 0x0a20
	13'h0511: q0 = 16'h3f00; // 0x0a22
	13'h0512: q0 = 16'h4247; // 0x0a24
	13'h0513: q0 = 16'h4246; // 0x0a26
	13'h0514: q0 = 16'h382e; // 0x0a28
	13'h0515: q0 = 16'h0008; // 0x0a2a
	13'h0516: q0 = 16'h362e; // 0x0a2c
	13'h0517: q0 = 16'h000a; // 0x0a2e
	13'h0518: q0 = 16'h4a44; // 0x0a30
	13'h0519: q0 = 16'h6c08; // 0x0a32
	13'h051a: q0 = 16'h7e01; // 0x0a34
	13'h051b: q0 = 16'h3004; // 0x0a36
	13'h051c: q0 = 16'h4440; // 0x0a38
	13'h051d: q0 = 16'h3800; // 0x0a3a
	13'h051e: q0 = 16'h4a43; // 0x0a3c
	13'h051f: q0 = 16'h6c08; // 0x0a3e
	13'h0520: q0 = 16'h7c01; // 0x0a40
	13'h0521: q0 = 16'h3003; // 0x0a42
	13'h0522: q0 = 16'h4440; // 0x0a44
	13'h0523: q0 = 16'h3600; // 0x0a46
	13'h0524: q0 = 16'hb87c; // 0x0a48
	13'h0525: q0 = 16'h000f; // 0x0a4a
	13'h0526: q0 = 16'h6e06; // 0x0a4c
	13'h0527: q0 = 16'hb67c; // 0x0a4e
	13'h0528: q0 = 16'h000f; // 0x0a50
	13'h0529: q0 = 16'h6f06; // 0x0a52
	13'h052a: q0 = 16'he244; // 0x0a54
	13'h052b: q0 = 16'he243; // 0x0a56
	13'h052c: q0 = 16'h60ee; // 0x0a58
	13'h052d: q0 = 16'h3004; // 0x0a5a
	13'h052e: q0 = 16'he940; // 0x0a5c
	13'h052f: q0 = 16'hd043; // 0x0a5e
	13'h0530: q0 = 16'h48c0; // 0x0a60
	13'h0531: q0 = 16'hd0bc; // 0x0a62
	13'h0532: q0 = 16'h0000; // 0x0a64
	13'h0533: q0 = 16'hc190; // 0x0a66
	13'h0534: q0 = 16'h2040; // 0x0a68
	13'h0535: q0 = 16'h1a10; // 0x0a6a
	13'h0536: q0 = 16'h4885; // 0x0a6c
	13'h0537: q0 = 16'h4a47; // 0x0a6e
	13'h0538: q0 = 16'h670a; // 0x0a70
	13'h0539: q0 = 16'h4a46; // 0x0a72
	13'h053a: q0 = 16'h6606; // 0x0a74
	13'h053b: q0 = 16'h7024; // 0x0a76
	13'h053c: q0 = 16'h9045; // 0x0a78
	13'h053d: q0 = 16'h3a00; // 0x0a7a
	13'h053e: q0 = 16'h4a46; // 0x0a7c
	13'h053f: q0 = 16'h670a; // 0x0a7e
	13'h0540: q0 = 16'h4a47; // 0x0a80
	13'h0541: q0 = 16'h6606; // 0x0a82
	13'h0542: q0 = 16'h7048; // 0x0a84
	13'h0543: q0 = 16'h9045; // 0x0a86
	13'h0544: q0 = 16'h3a00; // 0x0a88
	13'h0545: q0 = 16'h4a47; // 0x0a8a
	13'h0546: q0 = 16'h6708; // 0x0a8c
	13'h0547: q0 = 16'h4a46; // 0x0a8e
	13'h0548: q0 = 16'h6704; // 0x0a90
	13'h0549: q0 = 16'hda7c; // 0x0a92
	13'h054a: q0 = 16'h0024; // 0x0a94
	13'h054b: q0 = 16'hba7c; // 0x0a96
	13'h054c: q0 = 16'h0048; // 0x0a98
	13'h054d: q0 = 16'h6602; // 0x0a9a
	13'h054e: q0 = 16'h4245; // 0x0a9c
	13'h054f: q0 = 16'h3005; // 0x0a9e
	13'h0550: q0 = 16'h4a9f; // 0x0aa0
	13'h0551: q0 = 16'h4cdf; // 0x0aa2
	13'h0552: q0 = 16'h00f8; // 0x0aa4
	13'h0553: q0 = 16'h4e5e; // 0x0aa6
	13'h0554: q0 = 16'h4e75; // 0x0aa8
	13'h0555: q0 = 16'h4e56; // 0x0aaa
	13'h0556: q0 = 16'hfff6; // 0x0aac
	13'h0557: q0 = 16'h48e7; // 0x0aae
	13'h0558: q0 = 16'h1f1c; // 0x0ab0
	13'h0559: q0 = 16'h422e; // 0x0ab2
	13'h055a: q0 = 16'hfff6; // 0x0ab4
	13'h055b: q0 = 16'h4244; // 0x0ab6
	13'h055c: q0 = 16'h287c; // 0x0ab8
	13'h055d: q0 = 16'h0001; // 0x0aba
	13'h055e: q0 = 16'h87e0; // 0x0abc
	13'h055f: q0 = 16'h267c; // 0x0abe
	13'h0560: q0 = 16'h0001; // 0x0ac0
	13'h0561: q0 = 16'h892a; // 0x0ac2
	13'h0562: q0 = 16'hb87c; // 0x0ac4
	13'h0563: q0 = 16'h0005; // 0x0ac6
	13'h0564: q0 = 16'h6c28; // 0x0ac8
	13'h0565: q0 = 16'h3e84; // 0x0aca
	13'h0566: q0 = 16'h0657; // 0x0acc
	13'h0567: q0 = 16'h0029; // 0x0ace
	13'h0568: q0 = 16'h2f0c; // 0x0ad0
	13'h0569: q0 = 16'h4eb9; // 0x0ad2
	13'h056a: q0 = 16'h0000; // 0x0ad4
	13'h056b: q0 = 16'h78f6; // 0x0ad6
	13'h056c: q0 = 16'h4a9f; // 0x0ad8
	13'h056d: q0 = 16'hb87c; // 0x0ada
	13'h056e: q0 = 16'h0003; // 0x0adc
	13'h056f: q0 = 16'h6c06; // 0x0ade
	13'h0570: q0 = 16'h41ee; // 0x0ae0
	13'h0571: q0 = 16'hfff6; // 0x0ae2
	13'h0572: q0 = 16'h2688; // 0x0ae4
	13'h0573: q0 = 16'h5244; // 0x0ae6
	13'h0574: q0 = 16'hd9fc; // 0x0ae8
	13'h0575: q0 = 16'h0000; // 0x0aea
	13'h0576: q0 = 16'h0020; // 0x0aec
	13'h0577: q0 = 16'h588b; // 0x0aee
	13'h0578: q0 = 16'h60d2; // 0x0af0
	13'h0579: q0 = 16'h2a7c; // 0x0af2
	13'h057a: q0 = 16'h0001; // 0x0af4
	13'h057b: q0 = 16'h7f2c; // 0x0af6
	13'h057c: q0 = 16'h4279; // 0x0af8
	13'h057d: q0 = 16'h0001; // 0x0afa
	13'h057e: q0 = 16'h8054; // 0x0afc
	13'h057f: q0 = 16'h23fc; // 0x0afe
	13'h0580: q0 = 16'h0001; // 0x0b00
	13'h0581: q0 = 16'h8628; // 0x0b02
	13'h0582: q0 = 16'h0001; // 0x0b04
	13'h0583: q0 = 16'h7fb8; // 0x0b06
	13'h0584: q0 = 16'h33f9; // 0x0b08
	13'h0585: q0 = 16'h0001; // 0x0b0a
	13'h0586: q0 = 16'h757a; // 0x0b0c
	13'h0587: q0 = 16'h0001; // 0x0b0e
	13'h0588: q0 = 16'h862a; // 0x0b10
	13'h0589: q0 = 16'h33ee; // 0x0b12
	13'h058a: q0 = 16'h0008; // 0x0b14
	13'h058b: q0 = 16'h0001; // 0x0b16
	13'h058c: q0 = 16'h8628; // 0x0b18
	13'h058d: q0 = 16'h4eb9; // 0x0b1a
	13'h058e: q0 = 16'h0000; // 0x0b1c
	13'h058f: q0 = 16'h0226; // 0x0b1e
	13'h0590: q0 = 16'h4eb9; // 0x0b20
	13'h0591: q0 = 16'h0000; // 0x0b22
	13'h0592: q0 = 16'hb3c6; // 0x0b24
	13'h0593: q0 = 16'h4eb9; // 0x0b26
	13'h0594: q0 = 16'h0000; // 0x0b28
	13'h0595: q0 = 16'h90d4; // 0x0b2a
	13'h0596: q0 = 16'h4eb9; // 0x0b2c
	13'h0597: q0 = 16'h0000; // 0x0b2e
	13'h0598: q0 = 16'h0ea2; // 0x0b30
	13'h0599: q0 = 16'h4eb9; // 0x0b32
	13'h059a: q0 = 16'h0000; // 0x0b34
	13'h059b: q0 = 16'h41ae; // 0x0b36
	13'h059c: q0 = 16'h4eb9; // 0x0b38
	13'h059d: q0 = 16'h0000; // 0x0b3a
	13'h059e: q0 = 16'h4754; // 0x0b3c
	13'h059f: q0 = 16'h4eb9; // 0x0b3e
	13'h05a0: q0 = 16'h0000; // 0x0b40
	13'h05a1: q0 = 16'h4dee; // 0x0b42
	13'h05a2: q0 = 16'h4eb9; // 0x0b44
	13'h05a3: q0 = 16'h0000; // 0x0b46
	13'h05a4: q0 = 16'h8330; // 0x0b48
	13'h05a5: q0 = 16'h4eb9; // 0x0b4a
	13'h05a6: q0 = 16'h0000; // 0x0b4c
	13'h05a7: q0 = 16'h5a9c; // 0x0b4e
	13'h05a8: q0 = 16'h4eb9; // 0x0b50
	13'h05a9: q0 = 16'h0000; // 0x0b52
	13'h05aa: q0 = 16'h2cba; // 0x0b54
	13'h05ab: q0 = 16'h4279; // 0x0b56
	13'h05ac: q0 = 16'h0001; // 0x0b58
	13'h05ad: q0 = 16'h7b9e; // 0x0b5a
	13'h05ae: q0 = 16'h4247; // 0x0b5c
	13'h05af: q0 = 16'h4a79; // 0x0b5e
	13'h05b0: q0 = 16'h0001; // 0x0b60
	13'h05b1: q0 = 16'h7f5e; // 0x0b62
	13'h05b2: q0 = 16'h664c; // 0x0b64
	13'h05b3: q0 = 16'h200e; // 0x0b66
	13'h05b4: q0 = 16'hd0bc; // 0x0b68
	13'h05b5: q0 = 16'hffff; // 0x0b6a
	13'h05b6: q0 = 16'hfffc; // 0x0b6c
	13'h05b7: q0 = 16'h2e80; // 0x0b6e
	13'h05b8: q0 = 16'h200e; // 0x0b70
	13'h05b9: q0 = 16'hd0bc; // 0x0b72
	13'h05ba: q0 = 16'hffff; // 0x0b74
	13'h05bb: q0 = 16'hfffe; // 0x0b76
	13'h05bc: q0 = 16'h2f00; // 0x0b78
	13'h05bd: q0 = 16'h4eb9; // 0x0b7a
	13'h05be: q0 = 16'h0000; // 0x0b7c
	13'h05bf: q0 = 16'h182a; // 0x0b7e
	13'h05c0: q0 = 16'h4a9f; // 0x0b80
	13'h05c1: q0 = 16'h4a40; // 0x0b82
	13'h05c2: q0 = 16'h662c; // 0x0b84
	13'h05c3: q0 = 16'h23fc; // 0x0b86
	13'h05c4: q0 = 16'h0000; // 0x0b88
	13'h05c5: q0 = 16'h0002; // 0x0b8a
	13'h05c6: q0 = 16'h0001; // 0x0b8c
	13'h05c7: q0 = 16'h7fc2; // 0x0b8e
	13'h05c8: q0 = 16'h4eb9; // 0x0b90
	13'h05c9: q0 = 16'h0000; // 0x0b92
	13'h05ca: q0 = 16'h18d0; // 0x0b94
	13'h05cb: q0 = 16'h4eb9; // 0x0b96
	13'h05cc: q0 = 16'h0000; // 0x0b98
	13'h05cd: q0 = 16'h12ba; // 0x0b9a
	13'h05ce: q0 = 16'h4ab9; // 0x0b9c
	13'h05cf: q0 = 16'h0001; // 0x0b9e
	13'h05d0: q0 = 16'h7fc2; // 0x0ba0
	13'h05d1: q0 = 16'h670c; // 0x0ba2
	13'h05d2: q0 = 16'h4a79; // 0x0ba4
	13'h05d3: q0 = 16'h0001; // 0x0ba6
	13'h05d4: q0 = 16'h7f5e; // 0x0ba8
	13'h05d5: q0 = 16'h6600; // 0x0baa
	13'h05d6: q0 = 16'h01c6; // 0x0bac
	13'h05d7: q0 = 16'h60ec; // 0x0bae
	13'h05d8: q0 = 16'h60ac; // 0x0bb0
	13'h05d9: q0 = 16'h4a79; // 0x0bb2
	13'h05da: q0 = 16'h0001; // 0x0bb4
	13'h05db: q0 = 16'h7f5e; // 0x0bb6
	13'h05dc: q0 = 16'h6600; // 0x0bb8
	13'h05dd: q0 = 16'h01b8; // 0x0bba
	13'h05de: q0 = 16'h23fc; // 0x0bbc
	13'h05df: q0 = 16'h0000; // 0x0bbe
	13'h05e0: q0 = 16'h0002; // 0x0bc0
	13'h05e1: q0 = 16'h0001; // 0x0bc2
	13'h05e2: q0 = 16'h7fc2; // 0x0bc4
	13'h05e3: q0 = 16'h33fc; // 0x0bc6
	13'h05e4: q0 = 16'h0001; // 0x0bc8
	13'h05e5: q0 = 16'h0001; // 0x0bca
	13'h05e6: q0 = 16'h805a; // 0x0bcc
	13'h05e7: q0 = 16'h3c39; // 0x0bce
	13'h05e8: q0 = 16'h0001; // 0x0bd0
	13'h05e9: q0 = 16'h8936; // 0x0bd2
	13'h05ea: q0 = 16'h3a39; // 0x0bd4
	13'h05eb: q0 = 16'h0001; // 0x0bd6
	13'h05ec: q0 = 16'h8938; // 0x0bd8
	13'h05ed: q0 = 16'h33fc; // 0x0bda
	13'h05ee: q0 = 16'h0001; // 0x0bdc
	13'h05ef: q0 = 16'h0001; // 0x0bde
	13'h05f0: q0 = 16'h8880; // 0x0be0
	13'h05f1: q0 = 16'h33fc; // 0x0be2
	13'h05f2: q0 = 16'h0001; // 0x0be4
	13'h05f3: q0 = 16'h0001; // 0x0be6
	13'h05f4: q0 = 16'h81fa; // 0x0be8
	13'h05f5: q0 = 16'h4a47; // 0x0bea
	13'h05f6: q0 = 16'h6600; // 0x0bec
	13'h05f7: q0 = 16'h0084; // 0x0bee
	13'h05f8: q0 = 16'h4257; // 0x0bf0
	13'h05f9: q0 = 16'h206d; // 0x0bf2
	13'h05fa: q0 = 16'h0024; // 0x0bf4
	13'h05fb: q0 = 16'h3f28; // 0x0bf6
	13'h05fc: q0 = 16'h0002; // 0x0bf8
	13'h05fd: q0 = 16'h206d; // 0x0bfa
	13'h05fe: q0 = 16'h0024; // 0x0bfc
	13'h05ff: q0 = 16'h3f10; // 0x0bfe
	13'h0600: q0 = 16'h4eb9; // 0x0c00
	13'h0601: q0 = 16'h0000; // 0x0c02
	13'h0602: q0 = 16'h8744; // 0x0c04
	13'h0603: q0 = 16'h4a9f; // 0x0c06
	13'h0604: q0 = 16'h4a40; // 0x0c08
	13'h0605: q0 = 16'h6634; // 0x0c0a
	13'h0606: q0 = 16'h200e; // 0x0c0c
	13'h0607: q0 = 16'hd0bc; // 0x0c0e
	13'h0608: q0 = 16'hffff; // 0x0c10
	13'h0609: q0 = 16'hfffc; // 0x0c12
	13'h060a: q0 = 16'h2e80; // 0x0c14
	13'h060b: q0 = 16'h200e; // 0x0c16
	13'h060c: q0 = 16'hd0bc; // 0x0c18
	13'h060d: q0 = 16'hffff; // 0x0c1a
	13'h060e: q0 = 16'hfffe; // 0x0c1c
	13'h060f: q0 = 16'h2f00; // 0x0c1e
	13'h0610: q0 = 16'h4eb9; // 0x0c20
	13'h0611: q0 = 16'h0000; // 0x0c22
	13'h0612: q0 = 16'h86be; // 0x0c24
	13'h0613: q0 = 16'h4a9f; // 0x0c26
	13'h0614: q0 = 16'h4a40; // 0x0c28
	13'h0615: q0 = 16'h6710; // 0x0c2a
	13'h0616: q0 = 16'h3c2e; // 0x0c2c
	13'h0617: q0 = 16'hfffe; // 0x0c2e
	13'h0618: q0 = 16'h3a2e; // 0x0c30
	13'h0619: q0 = 16'hfffc; // 0x0c32
	13'h061a: q0 = 16'h4279; // 0x0c34
	13'h061b: q0 = 16'h0001; // 0x0c36
	13'h061c: q0 = 16'h81fa; // 0x0c38
	13'h061d: q0 = 16'h6002; // 0x0c3a
	13'h061e: q0 = 16'h7e01; // 0x0c3c
	13'h061f: q0 = 16'h6032; // 0x0c3e
	13'h0620: q0 = 16'h200e; // 0x0c40
	13'h0621: q0 = 16'hd0bc; // 0x0c42
	13'h0622: q0 = 16'hffff; // 0x0c44
	13'h0623: q0 = 16'hfffc; // 0x0c46
	13'h0624: q0 = 16'h2e80; // 0x0c48
	13'h0625: q0 = 16'h200e; // 0x0c4a
	13'h0626: q0 = 16'hd0bc; // 0x0c4c
	13'h0627: q0 = 16'hffff; // 0x0c4e
	13'h0628: q0 = 16'hfffe; // 0x0c50
	13'h0629: q0 = 16'h2f00; // 0x0c52
	13'h062a: q0 = 16'h4eb9; // 0x0c54
	13'h062b: q0 = 16'h0000; // 0x0c56
	13'h062c: q0 = 16'h182a; // 0x0c58
	13'h062d: q0 = 16'h4a9f; // 0x0c5a
	13'h062e: q0 = 16'h4a40; // 0x0c5c
	13'h062f: q0 = 16'h6710; // 0x0c5e
	13'h0630: q0 = 16'h3c2e; // 0x0c60
	13'h0631: q0 = 16'hfffe; // 0x0c62
	13'h0632: q0 = 16'h3a2e; // 0x0c64
	13'h0633: q0 = 16'hfffc; // 0x0c66
	13'h0634: q0 = 16'h4279; // 0x0c68
	13'h0635: q0 = 16'h0001; // 0x0c6a
	13'h0636: q0 = 16'h8880; // 0x0c6c
	13'h0637: q0 = 16'h6002; // 0x0c6e
	13'h0638: q0 = 16'h7e01; // 0x0c70
	13'h0639: q0 = 16'h3e85; // 0x0c72
	13'h063a: q0 = 16'h206d; // 0x0c74
	13'h063b: q0 = 16'h0024; // 0x0c76
	13'h063c: q0 = 16'h3028; // 0x0c78
	13'h063d: q0 = 16'h0002; // 0x0c7a
	13'h063e: q0 = 16'h9157; // 0x0c7c
	13'h063f: q0 = 16'h3f06; // 0x0c7e
	13'h0640: q0 = 16'h206d; // 0x0c80
	13'h0641: q0 = 16'h0024; // 0x0c82
	13'h0642: q0 = 16'h3010; // 0x0c84
	13'h0643: q0 = 16'h9157; // 0x0c86
	13'h0644: q0 = 16'h4eb9; // 0x0c88
	13'h0645: q0 = 16'h0000; // 0x0c8a
	13'h0646: q0 = 16'h0a1c; // 0x0c8c
	13'h0647: q0 = 16'h4a5f; // 0x0c8e
	13'h0648: q0 = 16'h33c0; // 0x0c90
	13'h0649: q0 = 16'h0001; // 0x0c92
	13'h064a: q0 = 16'h8682; // 0x0c94
	13'h064b: q0 = 16'h4a79; // 0x0c96
	13'h064c: q0 = 16'h0001; // 0x0c98
	13'h064d: q0 = 16'h7f5e; // 0x0c9a
	13'h064e: q0 = 16'h6600; // 0x0c9c
	13'h064f: q0 = 16'h00d4; // 0x0c9e
	13'h0650: q0 = 16'h2d79; // 0x0ca0
	13'h0651: q0 = 16'h0000; // 0x0ca2
	13'h0652: q0 = 16'hc2e4; // 0x0ca4
	13'h0653: q0 = 16'hfff8; // 0x0ca6
	13'h0654: q0 = 16'h2039; // 0x0ca8
	13'h0655: q0 = 16'h0000; // 0x0caa
	13'h0656: q0 = 16'hc2e8; // 0x0cac
	13'h0657: q0 = 16'he380; // 0x0cae
	13'h0658: q0 = 16'h91ae; // 0x0cb0
	13'h0659: q0 = 16'hfff8; // 0x0cb2
	13'h065a: q0 = 16'h206e; // 0x0cb4
	13'h065b: q0 = 16'hfff8; // 0x0cb6
	13'h065c: q0 = 16'h3010; // 0x0cb8
	13'h065d: q0 = 16'he340; // 0x0cba
	13'h065e: q0 = 16'hb07c; // 0x0cbc
	13'h065f: q0 = 16'h5292; // 0x0cbe
	13'h0660: q0 = 16'h6708; // 0x0cc0
	13'h0661: q0 = 16'h33fc; // 0x0cc2
	13'h0662: q0 = 16'h0001; // 0x0cc4
	13'h0663: q0 = 16'h0001; // 0x0cc6
	13'h0664: q0 = 16'h77e8; // 0x0cc8
	13'h0665: q0 = 16'h4eb9; // 0x0cca
	13'h0666: q0 = 16'h0000; // 0x0ccc
	13'h0667: q0 = 16'h3434; // 0x0cce
	13'h0668: q0 = 16'h4eb9; // 0x0cd0
	13'h0669: q0 = 16'h0000; // 0x0cd2
	13'h066a: q0 = 16'h12ba; // 0x0cd4
	13'h066b: q0 = 16'h4eb9; // 0x0cd6
	13'h066c: q0 = 16'h0000; // 0x0cd8
	13'h066d: q0 = 16'h18d0; // 0x0cda
	13'h066e: q0 = 16'h4eb9; // 0x0cdc
	13'h066f: q0 = 16'h0000; // 0x0cde
	13'h0670: q0 = 16'h4820; // 0x0ce0
	13'h0671: q0 = 16'h4eb9; // 0x0ce2
	13'h0672: q0 = 16'h0000; // 0x0ce4
	13'h0673: q0 = 16'h909e; // 0x0ce6
	13'h0674: q0 = 16'h4eb9; // 0x0ce8
	13'h0675: q0 = 16'h0000; // 0x0cea
	13'h0676: q0 = 16'h3fcc; // 0x0cec
	13'h0677: q0 = 16'h4eb9; // 0x0cee
	13'h0678: q0 = 16'h0000; // 0x0cf0
	13'h0679: q0 = 16'h4738; // 0x0cf2
	13'h067a: q0 = 16'h4a40; // 0x0cf4
	13'h067b: q0 = 16'h6764; // 0x0cf6
	13'h067c: q0 = 16'h4eb9; // 0x0cf8
	13'h067d: q0 = 16'h0000; // 0x0cfa
	13'h067e: q0 = 16'h3396; // 0x0cfc
	13'h067f: q0 = 16'h4a40; // 0x0cfe
	13'h0680: q0 = 16'h675a; // 0x0d00
	13'h0681: q0 = 16'h4eb9; // 0x0d02
	13'h0682: q0 = 16'h0000; // 0x0d04
	13'h0683: q0 = 16'h16c2; // 0x0d06
	13'h0684: q0 = 16'h4a40; // 0x0d08
	13'h0685: q0 = 16'h6750; // 0x0d0a
	13'h0686: q0 = 16'h4eb9; // 0x0d0c
	13'h0687: q0 = 16'h0000; // 0x0d0e
	13'h0688: q0 = 16'h3fac; // 0x0d10
	13'h0689: q0 = 16'h4a40; // 0x0d12
	13'h068a: q0 = 16'h6746; // 0x0d14
	13'h068b: q0 = 16'h4eb9; // 0x0d16
	13'h068c: q0 = 16'h0000; // 0x0d18
	13'h068d: q0 = 16'h18d0; // 0x0d1a
	13'h068e: q0 = 16'h23f9; // 0x0d1c
	13'h068f: q0 = 16'h0000; // 0x0d1e
	13'h0690: q0 = 16'hc2ec; // 0x0d20
	13'h0691: q0 = 16'h0001; // 0x0d22
	13'h0692: q0 = 16'h7f60; // 0x0d24
	13'h0693: q0 = 16'h4ab9; // 0x0d26
	13'h0694: q0 = 16'h0001; // 0x0d28
	13'h0695: q0 = 16'h7f60; // 0x0d2a
	13'h0696: q0 = 16'h672c; // 0x0d2c
	13'h0697: q0 = 16'h23fc; // 0x0d2e
	13'h0698: q0 = 16'h0000; // 0x0d30
	13'h0699: q0 = 16'h0002; // 0x0d32
	13'h069a: q0 = 16'h0001; // 0x0d34
	13'h069b: q0 = 16'h7fc2; // 0x0d36
	13'h069c: q0 = 16'h4a79; // 0x0d38
	13'h069d: q0 = 16'h0001; // 0x0d3a
	13'h069e: q0 = 16'h7f5e; // 0x0d3c
	13'h069f: q0 = 16'h6632; // 0x0d3e
	13'h06a0: q0 = 16'h4eb9; // 0x0d40
	13'h06a1: q0 = 16'h0000; // 0x0d42
	13'h06a2: q0 = 16'h12ba; // 0x0d44
	13'h06a3: q0 = 16'h4ab9; // 0x0d46
	13'h06a4: q0 = 16'h0001; // 0x0d48
	13'h06a5: q0 = 16'h7fc2; // 0x0d4a
	13'h06a6: q0 = 16'h670a; // 0x0d4c
	13'h06a7: q0 = 16'h4a79; // 0x0d4e
	13'h06a8: q0 = 16'h0001; // 0x0d50
	13'h06a9: q0 = 16'h7f5e; // 0x0d52
	13'h06aa: q0 = 16'h661c; // 0x0d54
	13'h06ab: q0 = 16'h60ee; // 0x0d56
	13'h06ac: q0 = 16'h60cc; // 0x0d58
	13'h06ad: q0 = 16'h6016; // 0x0d5a
	13'h06ae: q0 = 16'h4ab9; // 0x0d5c
	13'h06af: q0 = 16'h0001; // 0x0d5e
	13'h06b0: q0 = 16'h7fc2; // 0x0d60
	13'h06b1: q0 = 16'h670a; // 0x0d62
	13'h06b2: q0 = 16'h4a79; // 0x0d64
	13'h06b3: q0 = 16'h0001; // 0x0d66
	13'h06b4: q0 = 16'h7f5e; // 0x0d68
	13'h06b5: q0 = 16'h6606; // 0x0d6a
	13'h06b6: q0 = 16'h60ee; // 0x0d6c
	13'h06b7: q0 = 16'h6000; // 0x0d6e
	13'h06b8: q0 = 16'hfe42; // 0x0d70
	13'h06b9: q0 = 16'h4a9f; // 0x0d72
	13'h06ba: q0 = 16'h4cdf; // 0x0d74
	13'h06bb: q0 = 16'h38f0; // 0x0d76
	13'h06bc: q0 = 16'h4e5e; // 0x0d78
	13'h06bd: q0 = 16'h4e75; // 0x0d7a
	13'h06be: q0 = 16'h4e56; // 0x0d7c
	13'h06bf: q0 = 16'hfffc; // 0x0d7e
	13'h06c0: q0 = 16'h2079; // 0x0d80
	13'h06c1: q0 = 16'h0001; // 0x0d82
	13'h06c2: q0 = 16'h7fb8; // 0x0d84
	13'h06c3: q0 = 16'h5268; // 0x0d86
	13'h06c4: q0 = 16'h0002; // 0x0d88
	13'h06c5: q0 = 16'h3ebc; // 0x0d8a
	13'h06c6: q0 = 16'h000b; // 0x0d8c
	13'h06c7: q0 = 16'h4eb9; // 0x0d8e
	13'h06c8: q0 = 16'h0000; // 0x0d90
	13'h06c9: q0 = 16'h549c; // 0x0d92
	13'h06ca: q0 = 16'h3039; // 0x0d94
	13'h06cb: q0 = 16'h0001; // 0x0d96
	13'h06cc: q0 = 16'h8054; // 0x0d98
	13'h06cd: q0 = 16'he340; // 0x0d9a
	13'h06ce: q0 = 16'h48c0; // 0x0d9c
	13'h06cf: q0 = 16'hd0bc; // 0x0d9e
	13'h06d0: q0 = 16'h0001; // 0x0da0
	13'h06d1: q0 = 16'h75da; // 0x0da2
	13'h06d2: q0 = 16'h2040; // 0x0da4
	13'h06d3: q0 = 16'h5250; // 0x0da6
	13'h06d4: q0 = 16'h2ebc; // 0x0da8
	13'h06d5: q0 = 16'h0000; // 0x0daa
	13'h06d6: q0 = 16'hc392; // 0x0dac
	13'h06d7: q0 = 16'h4eb9; // 0x0dae
	13'h06d8: q0 = 16'h0000; // 0x0db0
	13'h06d9: q0 = 16'h7ff8; // 0x0db2
	13'h06da: q0 = 16'h4e5e; // 0x0db4
	13'h06db: q0 = 16'h4e75; // 0x0db6
	13'h06dc: q0 = 16'h4e56; // 0x0db8
	13'h06dd: q0 = 16'hfffc; // 0x0dba
	13'h06de: q0 = 16'h48e7; // 0x0dbc
	13'h06df: q0 = 16'h071c; // 0x0dbe
	13'h06e0: q0 = 16'h2679; // 0x0dc0
	13'h06e1: q0 = 16'h0001; // 0x0dc2
	13'h06e2: q0 = 16'h7fb8; // 0x0dc4
	13'h06e3: q0 = 16'h33fc; // 0x0dc6
	13'h06e4: q0 = 16'h0001; // 0x0dc8
	13'h06e5: q0 = 16'h0001; // 0x0dca
	13'h06e6: q0 = 16'h7bd6; // 0x0dcc
	13'h06e7: q0 = 16'h23fc; // 0x0dce
	13'h06e8: q0 = 16'h0000; // 0x0dd0
	13'h06e9: q0 = 16'h0002; // 0x0dd2
	13'h06ea: q0 = 16'h0001; // 0x0dd4
	13'h06eb: q0 = 16'h7fc2; // 0x0dd6
	13'h06ec: q0 = 16'h2a7c; // 0x0dd8
	13'h06ed: q0 = 16'h0001; // 0x0dda
	13'h06ee: q0 = 16'h893e; // 0x0ddc
	13'h06ef: q0 = 16'h4247; // 0x0dde
	13'h06f0: q0 = 16'hbe79; // 0x0de0
	13'h06f1: q0 = 16'h0001; // 0x0de2
	13'h06f2: q0 = 16'h7fa8; // 0x0de4
	13'h06f3: q0 = 16'h6c00; // 0x0de6
	13'h06f4: q0 = 16'h008c; // 0x0de8
	13'h06f5: q0 = 16'h4a6d; // 0x0dea
	13'h06f6: q0 = 16'h0006; // 0x0dec
	13'h06f7: q0 = 16'h6778; // 0x0dee
	13'h06f8: q0 = 16'h0c6d; // 0x0df0
	13'h06f9: q0 = 16'h0005; // 0x0df2
	13'h06fa: q0 = 16'h0004; // 0x0df4
	13'h06fb: q0 = 16'h6770; // 0x0df6
	13'h06fc: q0 = 16'h3ebc; // 0x0df8
	13'h06fd: q0 = 16'h0001; // 0x0dfa
	13'h06fe: q0 = 16'h3f2d; // 0x0dfc
	13'h06ff: q0 = 16'h000a; // 0x0dfe
	13'h0700: q0 = 16'h3f2d; // 0x0e00
	13'h0701: q0 = 16'h0008; // 0x0e02
	13'h0702: q0 = 16'h4eb9; // 0x0e04
	13'h0703: q0 = 16'h0000; // 0x0e06
	13'h0704: q0 = 16'h37e6; // 0x0e08
	13'h0705: q0 = 16'h4a9f; // 0x0e0a
	13'h0706: q0 = 16'h2840; // 0x0e0c
	13'h0707: q0 = 16'h200c; // 0x0e0e
	13'h0708: q0 = 16'h6762; // 0x0e10
	13'h0709: q0 = 16'h302b; // 0x0e12
	13'h070a: q0 = 16'h0014; // 0x0e14
	13'h070b: q0 = 16'h906d; // 0x0e16
	13'h070c: q0 = 16'h0008; // 0x0e18
	13'h070d: q0 = 16'h3d40; // 0x0e1a
	13'h070e: q0 = 16'hfffe; // 0x0e1c
	13'h070f: q0 = 16'h302b; // 0x0e1e
	13'h0710: q0 = 16'h0016; // 0x0e20
	13'h0711: q0 = 16'h906d; // 0x0e22
	13'h0712: q0 = 16'h000a; // 0x0e24
	13'h0713: q0 = 16'h3d40; // 0x0e26
	13'h0714: q0 = 16'hfffc; // 0x0e28
	13'h0715: q0 = 16'h3c3c; // 0x0e2a
	13'h0716: q0 = 16'h0400; // 0x0e2c
	13'h0717: q0 = 16'h200e; // 0x0e2e
	13'h0718: q0 = 16'hd0bc; // 0x0e30
	13'h0719: q0 = 16'hffff; // 0x0e32
	13'h071a: q0 = 16'hfffc; // 0x0e34
	13'h071b: q0 = 16'h2e80; // 0x0e36
	13'h071c: q0 = 16'h200e; // 0x0e38
	13'h071d: q0 = 16'hd0bc; // 0x0e3a
	13'h071e: q0 = 16'hffff; // 0x0e3c
	13'h071f: q0 = 16'hfffe; // 0x0e3e
	13'h0720: q0 = 16'h2f00; // 0x0e40
	13'h0721: q0 = 16'h3f06; // 0x0e42
	13'h0722: q0 = 16'h4eb9; // 0x0e44
	13'h0723: q0 = 16'h0000; // 0x0e46
	13'h0724: q0 = 16'h09bc; // 0x0e48
	13'h0725: q0 = 16'h5c4f; // 0x0e4a
	13'h0726: q0 = 16'h3eab; // 0x0e4c
	13'h0727: q0 = 16'h0016; // 0x0e4e
	13'h0728: q0 = 16'h3f2b; // 0x0e50
	13'h0729: q0 = 16'h0014; // 0x0e52
	13'h072a: q0 = 16'h3f2e; // 0x0e54
	13'h072b: q0 = 16'hfffc; // 0x0e56
	13'h072c: q0 = 16'h3f2e; // 0x0e58
	13'h072d: q0 = 16'hfffe; // 0x0e5a
	13'h072e: q0 = 16'h2f0c; // 0x0e5c
	13'h072f: q0 = 16'h4eb9; // 0x0e5e
	13'h0730: q0 = 16'h0000; // 0x0e60
	13'h0731: q0 = 16'h3988; // 0x0e62
	13'h0732: q0 = 16'hdefc; // 0x0e64
	13'h0733: q0 = 16'h000a; // 0x0e66
	13'h0734: q0 = 16'hdbfc; // 0x0e68
	13'h0735: q0 = 16'h0000; // 0x0e6a
	13'h0736: q0 = 16'h0010; // 0x0e6c
	13'h0737: q0 = 16'h5247; // 0x0e6e
	13'h0738: q0 = 16'h6000; // 0x0e70
	13'h0739: q0 = 16'hff6e; // 0x0e72
	13'h073a: q0 = 16'h4eb9; // 0x0e74
	13'h073b: q0 = 16'h0000; // 0x0e76
	13'h073c: q0 = 16'h2fb4; // 0x0e78
	13'h073d: q0 = 16'h4eb9; // 0x0e7a
	13'h073e: q0 = 16'h0000; // 0x0e7c
	13'h073f: q0 = 16'h3396; // 0x0e7e
	13'h0740: q0 = 16'h4a40; // 0x0e80
	13'h0741: q0 = 16'h660e; // 0x0e82
	13'h0742: q0 = 16'h4ab9; // 0x0e84
	13'h0743: q0 = 16'h0001; // 0x0e86
	13'h0744: q0 = 16'h7fc2; // 0x0e88
	13'h0745: q0 = 16'h6702; // 0x0e8a
	13'h0746: q0 = 16'h60f6; // 0x0e8c
	13'h0747: q0 = 16'h6000; // 0x0e8e
	13'h0748: q0 = 16'hff3e; // 0x0e90
	13'h0749: q0 = 16'h4279; // 0x0e92
	13'h074a: q0 = 16'h0001; // 0x0e94
	13'h074b: q0 = 16'h7bd6; // 0x0e96
	13'h074c: q0 = 16'h4a9f; // 0x0e98
	13'h074d: q0 = 16'h4cdf; // 0x0e9a
	13'h074e: q0 = 16'h38c0; // 0x0e9c
	13'h074f: q0 = 16'h4e5e; // 0x0e9e
	13'h0750: q0 = 16'h4e75; // 0x0ea0
	13'h0751: q0 = 16'h4e56; // 0x0ea2
	13'h0752: q0 = 16'hffdc; // 0x0ea4
	13'h0753: q0 = 16'h48e7; // 0x0ea6
	13'h0754: q0 = 16'h0f0c; // 0x0ea8
	13'h0755: q0 = 16'h422e; // 0x0eaa
	13'h0756: q0 = 16'hfffe; // 0x0eac
	13'h0757: q0 = 16'h4bee; // 0x0eae
	13'h0758: q0 = 16'hffde; // 0x0eb0
	13'h0759: q0 = 16'h49ee; // 0x0eb2
	13'h075a: q0 = 16'hfffd; // 0x0eb4
	13'h075b: q0 = 16'h7c05; // 0x0eb6
	13'h075c: q0 = 16'hbc7c; // 0x0eb8
	13'h075d: q0 = 16'h001e; // 0x0eba
	13'h075e: q0 = 16'h6e00; // 0x0ebc
	13'h075f: q0 = 16'h0098; // 0x0ebe
	13'h0760: q0 = 16'hbc7c; // 0x0ec0
	13'h0761: q0 = 16'h0005; // 0x0ec2
	13'h0762: q0 = 16'h6614; // 0x0ec4
	13'h0763: q0 = 16'h1abc; // 0x0ec6
	13'h0764: q0 = 16'h003e; // 0x0ec8
	13'h0765: q0 = 16'h18bc; // 0x0eca
	13'h0766: q0 = 16'h003c; // 0x0ecc
	13'h0767: q0 = 16'h1a3c; // 0x0ece
	13'h0768: q0 = 16'h001b; // 0x0ed0
	13'h0769: q0 = 16'h3d7c; // 0x0ed2
	13'h076a: q0 = 16'h0001; // 0x0ed4
	13'h076b: q0 = 16'hffdc; // 0x0ed6
	13'h076c: q0 = 16'h6038; // 0x0ed8
	13'h076d: q0 = 16'hbc7c; // 0x0eda
	13'h076e: q0 = 16'h001e; // 0x0edc
	13'h076f: q0 = 16'h6614; // 0x0ede
	13'h0770: q0 = 16'h1abc; // 0x0ee0
	13'h0771: q0 = 16'h003d; // 0x0ee2
	13'h0772: q0 = 16'h18bc; // 0x0ee4
	13'h0773: q0 = 16'h003b; // 0x0ee6
	13'h0774: q0 = 16'h1a3c; // 0x0ee8
	13'h0775: q0 = 16'h0018; // 0x0eea
	13'h0776: q0 = 16'h3d7c; // 0x0eec
	13'h0777: q0 = 16'h0001; // 0x0eee
	13'h0778: q0 = 16'hffdc; // 0x0ef0
	13'h0779: q0 = 16'h601e; // 0x0ef2
	13'h077a: q0 = 16'hbc7c; // 0x0ef4
	13'h077b: q0 = 16'h0006; // 0x0ef6
	13'h077c: q0 = 16'h6614; // 0x0ef8
	13'h077d: q0 = 16'h1abc; // 0x0efa
	13'h077e: q0 = 16'h001a; // 0x0efc
	13'h077f: q0 = 16'h18bc; // 0x0efe
	13'h0780: q0 = 16'h0019; // 0x0f00
	13'h0781: q0 = 16'h1a3c; // 0x0f02
	13'h0782: q0 = 16'h0040; // 0x0f04
	13'h0783: q0 = 16'h3d7c; // 0x0f06
	13'h0784: q0 = 16'h0001; // 0x0f08
	13'h0785: q0 = 16'hffdc; // 0x0f0a
	13'h0786: q0 = 16'h6004; // 0x0f0c
	13'h0787: q0 = 16'h426e; // 0x0f0e
	13'h0788: q0 = 16'hffdc; // 0x0f10
	13'h0789: q0 = 16'h4a6e; // 0x0f12
	13'h078a: q0 = 16'hffdc; // 0x0f14
	13'h078b: q0 = 16'h671a; // 0x0f16
	13'h078c: q0 = 16'h7e01; // 0x0f18
	13'h078d: q0 = 16'hbe7c; // 0x0f1a
	13'h078e: q0 = 16'h001f; // 0x0f1c
	13'h078f: q0 = 16'h6c12; // 0x0f1e
	13'h0790: q0 = 16'h3207; // 0x0f20
	13'h0791: q0 = 16'h48c1; // 0x0f22
	13'h0792: q0 = 16'h200e; // 0x0f24
	13'h0793: q0 = 16'hd081; // 0x0f26
	13'h0794: q0 = 16'h2040; // 0x0f28
	13'h0795: q0 = 16'h1145; // 0x0f2a
	13'h0796: q0 = 16'hffde; // 0x0f2c
	13'h0797: q0 = 16'h5247; // 0x0f2e
	13'h0798: q0 = 16'h60e8; // 0x0f30
	13'h0799: q0 = 16'h3ebc; // 0x0f32
	13'h079a: q0 = 16'h0039; // 0x0f34
	13'h079b: q0 = 16'h4267; // 0x0f36
	13'h079c: q0 = 16'h4267; // 0x0f38
	13'h079d: q0 = 16'h3f06; // 0x0f3a
	13'h079e: q0 = 16'h200e; // 0x0f3c
	13'h079f: q0 = 16'hd0bc; // 0x0f3e
	13'h07a0: q0 = 16'hffff; // 0x0f40
	13'h07a1: q0 = 16'hffde; // 0x0f42
	13'h07a2: q0 = 16'h2f00; // 0x0f44
	13'h07a3: q0 = 16'h4eb9; // 0x0f46
	13'h07a4: q0 = 16'h0000; // 0x0f48
	13'h07a5: q0 = 16'h026c; // 0x0f4a
	13'h07a6: q0 = 16'hdefc; // 0x0f4c
	13'h07a7: q0 = 16'h000a; // 0x0f4e
	13'h07a8: q0 = 16'h5246; // 0x0f50
	13'h07a9: q0 = 16'h6000; // 0x0f52
	13'h07aa: q0 = 16'hff64; // 0x0f54
	13'h07ab: q0 = 16'h4a9f; // 0x0f56
	13'h07ac: q0 = 16'h4cdf; // 0x0f58
	13'h07ad: q0 = 16'h30e0; // 0x0f5a
	13'h07ae: q0 = 16'h4e5e; // 0x0f5c
	13'h07af: q0 = 16'h4e75; // 0x0f5e
	13'h07b0: q0 = 16'h4e56; // 0x0f60
	13'h07b1: q0 = 16'h0000; // 0x0f62
	13'h07b2: q0 = 16'h48e7; // 0x0f64
	13'h07b3: q0 = 16'h0f04; // 0x0f66
	13'h07b4: q0 = 16'h2a6e; // 0x0f68
	13'h07b5: q0 = 16'h0008; // 0x0f6a
	13'h07b6: q0 = 16'h3e2d; // 0x0f6c
	13'h07b7: q0 = 16'h0004; // 0x0f6e
	13'h07b8: q0 = 16'h3c2d; // 0x0f70
	13'h07b9: q0 = 16'h0006; // 0x0f72
	13'h07ba: q0 = 16'h3a15; // 0x0f74
	13'h07bb: q0 = 16'hbc7c; // 0x0f76
	13'h07bc: q0 = 16'h0001; // 0x0f78
	13'h07bd: q0 = 16'h6610; // 0x0f7a
	13'h07be: q0 = 16'hbe7c; // 0x0f7c
	13'h07bf: q0 = 16'h0002; // 0x0f7e
	13'h07c0: q0 = 16'h670a; // 0x0f80
	13'h07c1: q0 = 16'hbe7c; // 0x0f82
	13'h07c2: q0 = 16'h0001; // 0x0f84
	13'h07c3: q0 = 16'h6704; // 0x0f86
	13'h07c4: q0 = 16'h9a7c; // 0x0f88
	13'h07c5: q0 = 16'h0200; // 0x0f8a
	13'h07c6: q0 = 16'h3b45; // 0x0f8c
	13'h07c7: q0 = 16'h0008; // 0x0f8e
	13'h07c8: q0 = 16'h3a2d; // 0x0f90
	13'h07c9: q0 = 16'h0002; // 0x0f92
	13'h07ca: q0 = 16'hbc7c; // 0x0f94
	13'h07cb: q0 = 16'h0004; // 0x0f96
	13'h07cc: q0 = 16'h6e04; // 0x0f98
	13'h07cd: q0 = 16'h9a7c; // 0x0f9a
	13'h07ce: q0 = 16'h0200; // 0x0f9c
	13'h07cf: q0 = 16'h3b45; // 0x0f9e
	13'h07d0: q0 = 16'h000a; // 0x0fa0
	13'h07d1: q0 = 16'hbc7c; // 0x0fa2
	13'h07d2: q0 = 16'h0001; // 0x0fa4
	13'h07d3: q0 = 16'h6606; // 0x0fa6
	13'h07d4: q0 = 16'h3a3c; // 0x0fa8
	13'h07d5: q0 = 16'h0400; // 0x0faa
	13'h07d6: q0 = 16'h6004; // 0x0fac
	13'h07d7: q0 = 16'h3a3c; // 0x0fae
	13'h07d8: q0 = 16'h0600; // 0x0fb0
	13'h07d9: q0 = 16'h3b45; // 0x0fb2
	13'h07da: q0 = 16'h000c; // 0x0fb4
	13'h07db: q0 = 16'hbc7c; // 0x0fb6
	13'h07dc: q0 = 16'h0004; // 0x0fb8
	13'h07dd: q0 = 16'h6e06; // 0x0fba
	13'h07de: q0 = 16'h3a3c; // 0x0fbc
	13'h07df: q0 = 16'h0400; // 0x0fbe
	13'h07e0: q0 = 16'h6004; // 0x0fc0
	13'h07e1: q0 = 16'h3a3c; // 0x0fc2
	13'h07e2: q0 = 16'h0600; // 0x0fc4
	13'h07e3: q0 = 16'h3b45; // 0x0fc6
	13'h07e4: q0 = 16'h000e; // 0x0fc8
	13'h07e5: q0 = 16'h4a9f; // 0x0fca
	13'h07e6: q0 = 16'h4cdf; // 0x0fcc
	13'h07e7: q0 = 16'h20e0; // 0x0fce
	13'h07e8: q0 = 16'h4e5e; // 0x0fd0
	13'h07e9: q0 = 16'h4e75; // 0x0fd2
	13'h07ea: q0 = 16'h4e56; // 0x0fd4
	13'h07eb: q0 = 16'hfffc; // 0x0fd6
	13'h07ec: q0 = 16'h4279; // 0x0fd8
	13'h07ed: q0 = 16'h0001; // 0x0fda
	13'h07ee: q0 = 16'h893a; // 0x0fdc
	13'h07ef: q0 = 16'h4279; // 0x0fde
	13'h07f0: q0 = 16'h0001; // 0x0fe0
	13'h07f1: q0 = 16'h7bd8; // 0x0fe2
	13'h07f2: q0 = 16'h4279; // 0x0fe4
	13'h07f3: q0 = 16'h0001; // 0x0fe6
	13'h07f4: q0 = 16'h7594; // 0x0fe8
	13'h07f5: q0 = 16'h4279; // 0x0fea
	13'h07f6: q0 = 16'h0001; // 0x0fec
	13'h07f7: q0 = 16'h75e6; // 0x0fee
	13'h07f8: q0 = 16'h4240; // 0x0ff0
	13'h07f9: q0 = 16'h33c0; // 0x0ff2
	13'h07fa: q0 = 16'h0001; // 0x0ff4
	13'h07fb: q0 = 16'h8056; // 0x0ff6
	13'h07fc: q0 = 16'h33c0; // 0x0ff8
	13'h07fd: q0 = 16'h0001; // 0x0ffa
	13'h07fe: q0 = 16'h8620; // 0x0ffc
	13'h07ff: q0 = 16'h33c0; // 0x0ffe
	13'h0800: q0 = 16'h0001; // 0x1000
	13'h0801: q0 = 16'h85fa; // 0x1002
	13'h0802: q0 = 16'h4240; // 0x1004
	13'h0803: q0 = 16'h33c0; // 0x1006
	13'h0804: q0 = 16'h0001; // 0x1008
	13'h0805: q0 = 16'h81f2; // 0x100a
	13'h0806: q0 = 16'h33c0; // 0x100c
	13'h0807: q0 = 16'h0001; // 0x100e
	13'h0808: q0 = 16'h86ac; // 0x1010
	13'h0809: q0 = 16'h33c0; // 0x1012
	13'h080a: q0 = 16'h0001; // 0x1014
	13'h080b: q0 = 16'h8674; // 0x1016
	13'h080c: q0 = 16'h4240; // 0x1018
	13'h080d: q0 = 16'h33c0; // 0x101a
	13'h080e: q0 = 16'h0001; // 0x101c
	13'h080f: q0 = 16'h867c; // 0x101e
	13'h0810: q0 = 16'h33c0; // 0x1020
	13'h0811: q0 = 16'h0001; // 0x1022
	13'h0812: q0 = 16'h861a; // 0x1024
	13'h0813: q0 = 16'h4e5e; // 0x1026
	13'h0814: q0 = 16'h4e75; // 0x1028
	13'h0815: q0 = 16'h4e56; // 0x102a
	13'h0816: q0 = 16'hfff0; // 0x102c
	13'h0817: q0 = 16'h48e7; // 0x102e
	13'h0818: q0 = 16'h3f04; // 0x1030
	13'h0819: q0 = 16'h4a79; // 0x1032
	13'h081a: q0 = 16'h0001; // 0x1034
	13'h081b: q0 = 16'h8a7c; // 0x1036
	13'h081c: q0 = 16'h6706; // 0x1038
	13'h081d: q0 = 16'h4eb9; // 0x103a
	13'h081e: q0 = 16'h0000; // 0x103c
	13'h081f: q0 = 16'h9c8a; // 0x103e
	13'h0820: q0 = 16'h4244; // 0x1040
	13'h0821: q0 = 16'hb87c; // 0x1042
	13'h0822: q0 = 16'h0008; // 0x1044
	13'h0823: q0 = 16'h6c20; // 0x1046
	13'h0824: q0 = 16'h3004; // 0x1048
	13'h0825: q0 = 16'he340; // 0x104a
	13'h0826: q0 = 16'h48c0; // 0x104c
	13'h0827: q0 = 16'hd08e; // 0x104e
	13'h0828: q0 = 16'h2040; // 0x1050
	13'h0829: q0 = 16'h3204; // 0x1052
	13'h082a: q0 = 16'he341; // 0x1054
	13'h082b: q0 = 16'h48c1; // 0x1056
	13'h082c: q0 = 16'hd2bc; // 0x1058
	13'h082d: q0 = 16'h0001; // 0x105a
	13'h082e: q0 = 16'h805c; // 0x105c
	13'h082f: q0 = 16'h2241; // 0x105e
	13'h0830: q0 = 16'h3151; // 0x1060
	13'h0831: q0 = 16'hfff0; // 0x1062
	13'h0832: q0 = 16'h5244; // 0x1064
	13'h0833: q0 = 16'h60da; // 0x1066
	13'h0834: q0 = 16'h4a6e; // 0x1068
	13'h0835: q0 = 16'hfff0; // 0x106a
	13'h0836: q0 = 16'h6612; // 0x106c
	13'h0837: q0 = 16'h4a6e; // 0x106e
	13'h0838: q0 = 16'hfff2; // 0x1070
	13'h0839: q0 = 16'h670c; // 0x1072
	13'h083a: q0 = 16'h33fc; // 0x1074
	13'h083b: q0 = 16'h0002; // 0x1076
	13'h083c: q0 = 16'h0001; // 0x1078
	13'h083d: q0 = 16'h7594; // 0x107a
	13'h083e: q0 = 16'h6000; // 0x107c
	13'h083f: q0 = 16'h01de; // 0x107e
	13'h0840: q0 = 16'h2a79; // 0x1080
	13'h0841: q0 = 16'h0000; // 0x1082
	13'h0842: q0 = 16'hc552; // 0x1084
	13'h0843: q0 = 16'h3e15; // 0x1086
	13'h0844: q0 = 16'hce7c; // 0x1088
	13'h0845: q0 = 16'h0002; // 0x108a
	13'h0846: q0 = 16'h3c15; // 0x108c
	13'h0847: q0 = 16'hcc7c; // 0x108e
	13'h0848: q0 = 16'h0001; // 0x1090
	13'h0849: q0 = 16'h3a15; // 0x1092
	13'h084a: q0 = 16'hca7c; // 0x1094
	13'h084b: q0 = 16'h0010; // 0x1096
	13'h084c: q0 = 16'h4243; // 0x1098
	13'h084d: q0 = 16'hbe79; // 0x109a
	13'h084e: q0 = 16'h0001; // 0x109c
	13'h084f: q0 = 16'h8620; // 0x109e
	13'h0850: q0 = 16'h665a; // 0x10a0
	13'h0851: q0 = 16'h3039; // 0x10a2
	13'h0852: q0 = 16'h0001; // 0x10a4
	13'h0853: q0 = 16'h86ac; // 0x10a6
	13'h0854: q0 = 16'h3207; // 0x10a8
	13'h0855: q0 = 16'hb340; // 0x10aa
	13'h0856: q0 = 16'hc079; // 0x10ac
	13'h0857: q0 = 16'h0001; // 0x10ae
	13'h0858: q0 = 16'h86ac; // 0x10b0
	13'h0859: q0 = 16'h6742; // 0x10b2
	13'h085a: q0 = 16'h4a6e; // 0x10b4
	13'h085b: q0 = 16'hfff6; // 0x10b6
	13'h085c: q0 = 16'h660e; // 0x10b8
	13'h085d: q0 = 16'h4a6e; // 0x10ba
	13'h085e: q0 = 16'hfff4; // 0x10bc
	13'h085f: q0 = 16'h6604; // 0x10be
	13'h0860: q0 = 16'h7801; // 0x10c0
	13'h0861: q0 = 16'h6002; // 0x10c2
	13'h0862: q0 = 16'h7804; // 0x10c4
	13'h0863: q0 = 16'h600c; // 0x10c6
	13'h0864: q0 = 16'h4a6e; // 0x10c8
	13'h0865: q0 = 16'hfff4; // 0x10ca
	13'h0866: q0 = 16'h6604; // 0x10cc
	13'h0867: q0 = 16'h7805; // 0x10ce
	13'h0868: q0 = 16'h6002; // 0x10d0
	13'h0869: q0 = 16'h7806; // 0x10d2
	13'h086a: q0 = 16'hd644; // 0x10d4
	13'h086b: q0 = 16'h52b9; // 0x10d6
	13'h086c: q0 = 16'h0001; // 0x10d8
	13'h086d: q0 = 16'h75a2; // 0x10da
	13'h086e: q0 = 16'h33fc; // 0x10dc
	13'h086f: q0 = 16'h0004; // 0x10de
	13'h0870: q0 = 16'h0001; // 0x10e0
	13'h0871: q0 = 16'h867c; // 0x10e2
	13'h0872: q0 = 16'h0c79; // 0x10e4
	13'h0873: q0 = 16'h0001; // 0x10e6
	13'h0874: q0 = 16'h0001; // 0x10e8
	13'h0875: q0 = 16'h7592; // 0x10ea
	13'h0876: q0 = 16'h6608; // 0x10ec
	13'h0877: q0 = 16'h33fc; // 0x10ee
	13'h0878: q0 = 16'h0004; // 0x10f0
	13'h0879: q0 = 16'h0001; // 0x10f2
	13'h087a: q0 = 16'h861a; // 0x10f4
	13'h087b: q0 = 16'h33c7; // 0x10f6
	13'h087c: q0 = 16'h0001; // 0x10f8
	13'h087d: q0 = 16'h86ac; // 0x10fa
	13'h087e: q0 = 16'hbc79; // 0x10fc
	13'h087f: q0 = 16'h0001; // 0x10fe
	13'h0880: q0 = 16'h85fa; // 0x1100
	13'h0881: q0 = 16'h6640; // 0x1102
	13'h0882: q0 = 16'h3039; // 0x1104
	13'h0883: q0 = 16'h0001; // 0x1106
	13'h0884: q0 = 16'h8674; // 0x1108
	13'h0885: q0 = 16'h3206; // 0x110a
	13'h0886: q0 = 16'hb340; // 0x110c
	13'h0887: q0 = 16'hc079; // 0x110e
	13'h0888: q0 = 16'h0001; // 0x1110
	13'h0889: q0 = 16'h8674; // 0x1112
	13'h088a: q0 = 16'h6728; // 0x1114
	13'h088b: q0 = 16'h302e; // 0x1116
	13'h088c: q0 = 16'hfff8; // 0x1118
	13'h088d: q0 = 16'h5240; // 0x111a
	13'h088e: q0 = 16'hd640; // 0x111c
	13'h088f: q0 = 16'h52b9; // 0x111e
	13'h0890: q0 = 16'h0001; // 0x1120
	13'h0891: q0 = 16'h75a6; // 0x1122
	13'h0892: q0 = 16'h33fc; // 0x1124
	13'h0893: q0 = 16'h0004; // 0x1126
	13'h0894: q0 = 16'h0001; // 0x1128
	13'h0895: q0 = 16'h861a; // 0x112a
	13'h0896: q0 = 16'h0c79; // 0x112c
	13'h0897: q0 = 16'h0001; // 0x112e
	13'h0898: q0 = 16'h0001; // 0x1130
	13'h0899: q0 = 16'h7592; // 0x1132
	13'h089a: q0 = 16'h6608; // 0x1134
	13'h089b: q0 = 16'h33fc; // 0x1136
	13'h089c: q0 = 16'h0004; // 0x1138
	13'h089d: q0 = 16'h0001; // 0x113a
	13'h089e: q0 = 16'h867c; // 0x113c
	13'h089f: q0 = 16'h33c6; // 0x113e
	13'h08a0: q0 = 16'h0001; // 0x1140
	13'h08a1: q0 = 16'h8674; // 0x1142
	13'h08a2: q0 = 16'hba79; // 0x1144
	13'h08a3: q0 = 16'h0001; // 0x1146
	13'h08a4: q0 = 16'h8056; // 0x1148
	13'h08a5: q0 = 16'h663a; // 0x114a
	13'h08a6: q0 = 16'h3039; // 0x114c
	13'h08a7: q0 = 16'h0001; // 0x114e
	13'h08a8: q0 = 16'h81f2; // 0x1150
	13'h08a9: q0 = 16'h3205; // 0x1152
	13'h08aa: q0 = 16'hb340; // 0x1154
	13'h08ab: q0 = 16'hc079; // 0x1156
	13'h08ac: q0 = 16'h0001; // 0x1158
	13'h08ad: q0 = 16'h81f2; // 0x115a
	13'h08ae: q0 = 16'h671e; // 0x115c
	13'h08af: q0 = 16'h5279; // 0x115e
	13'h08b0: q0 = 16'h0001; // 0x1160
	13'h08b1: q0 = 16'h7594; // 0x1162
	13'h08b2: q0 = 16'h52b9; // 0x1164
	13'h08b3: q0 = 16'h0001; // 0x1166
	13'h08b4: q0 = 16'h75ae; // 0x1168
	13'h08b5: q0 = 16'h52b9; // 0x116a
	13'h08b6: q0 = 16'h0001; // 0x116c
	13'h08b7: q0 = 16'h75ce; // 0x116e
	13'h08b8: q0 = 16'h2ebc; // 0x1170
	13'h08b9: q0 = 16'h0000; // 0x1172
	13'h08ba: q0 = 16'hc53a; // 0x1174
	13'h08bb: q0 = 16'h4eb9; // 0x1176
	13'h08bc: q0 = 16'h0000; // 0x1178
	13'h08bd: q0 = 16'h7e06; // 0x117a
	13'h08be: q0 = 16'h33f9; // 0x117c
	13'h08bf: q0 = 16'h0001; // 0x117e
	13'h08c0: q0 = 16'h8056; // 0x1180
	13'h08c1: q0 = 16'h0001; // 0x1182
	13'h08c2: q0 = 16'h81f2; // 0x1184
	13'h08c3: q0 = 16'h33c6; // 0x1186
	13'h08c4: q0 = 16'h0001; // 0x1188
	13'h08c5: q0 = 16'h85fa; // 0x118a
	13'h08c6: q0 = 16'h33c7; // 0x118c
	13'h08c7: q0 = 16'h0001; // 0x118e
	13'h08c8: q0 = 16'h8620; // 0x1190
	13'h08c9: q0 = 16'h33c5; // 0x1192
	13'h08ca: q0 = 16'h0001; // 0x1194
	13'h08cb: q0 = 16'h8056; // 0x1196
	13'h08cc: q0 = 16'hd779; // 0x1198
	13'h08cd: q0 = 16'h0001; // 0x119a
	13'h08ce: q0 = 16'h7bd8; // 0x119c
	13'h08cf: q0 = 16'hd779; // 0x119e
	13'h08d0: q0 = 16'h0001; // 0x11a0
	13'h08d1: q0 = 16'h893a; // 0x11a2
	13'h08d2: q0 = 16'h3c39; // 0x11a4
	13'h08d3: q0 = 16'h0001; // 0x11a6
	13'h08d4: q0 = 16'h893a; // 0x11a8
	13'h08d5: q0 = 16'h3e39; // 0x11aa
	13'h08d6: q0 = 16'h0001; // 0x11ac
	13'h08d7: q0 = 16'h7bd8; // 0x11ae
	13'h08d8: q0 = 16'h302e; // 0x11b0
	13'h08d9: q0 = 16'hfffc; // 0x11b2
	13'h08da: q0 = 16'hb06e; // 0x11b4
	13'h08db: q0 = 16'hfffe; // 0x11b6
	13'h08dc: q0 = 16'h6730; // 0x11b8
	13'h08dd: q0 = 16'h4a6e; // 0x11ba
	13'h08de: q0 = 16'hfffc; // 0x11bc
	13'h08df: q0 = 16'h6714; // 0x11be
	13'h08e0: q0 = 16'hbe7c; // 0x11c0
	13'h08e1: q0 = 16'h0004; // 0x11c2
	13'h08e2: q0 = 16'h6d0c; // 0x11c4
	13'h08e3: q0 = 16'h302e; // 0x11c6
	13'h08e4: q0 = 16'hfffa; // 0x11c8
	13'h08e5: q0 = 16'h5240; // 0x11ca
	13'h08e6: q0 = 16'hdc40; // 0x11cc
	13'h08e7: q0 = 16'h5947; // 0x11ce
	13'h08e8: q0 = 16'h60ee; // 0x11d0
	13'h08e9: q0 = 16'h6016; // 0x11d2
	13'h08ea: q0 = 16'h4a6e; // 0x11d4
	13'h08eb: q0 = 16'hfffa; // 0x11d6
	13'h08ec: q0 = 16'h6704; // 0x11d8
	13'h08ed: q0 = 16'h7802; // 0x11da
	13'h08ee: q0 = 16'h6002; // 0x11dc
	13'h08ef: q0 = 16'h7805; // 0x11de
	13'h08f0: q0 = 16'hbe44; // 0x11e0
	13'h08f1: q0 = 16'h6d06; // 0x11e2
	13'h08f2: q0 = 16'h5246; // 0x11e4
	13'h08f3: q0 = 16'h9e44; // 0x11e6
	13'h08f4: q0 = 16'h60f6; // 0x11e8
	13'h08f5: q0 = 16'h4243; // 0x11ea
	13'h08f6: q0 = 16'h4a46; // 0x11ec
	13'h08f7: q0 = 16'h6f24; // 0x11ee
	13'h08f8: q0 = 16'h4a6e; // 0x11f0
	13'h08f9: q0 = 16'hfff0; // 0x11f2
	13'h08fa: q0 = 16'h6712; // 0x11f4
	13'h08fb: q0 = 16'h4a6e; // 0x11f6
	13'h08fc: q0 = 16'hfff2; // 0x11f8
	13'h08fd: q0 = 16'h660c; // 0x11fa
	13'h08fe: q0 = 16'hbc7c; // 0x11fc
	13'h08ff: q0 = 16'h0001; // 0x11fe
	13'h0900: q0 = 16'h6712; // 0x1200
	13'h0901: q0 = 16'h5243; // 0x1202
	13'h0902: q0 = 16'h5546; // 0x1204
	13'h0903: q0 = 16'h600a; // 0x1206
	13'h0904: q0 = 16'h5346; // 0x1208
	13'h0905: q0 = 16'h302e; // 0x120a
	13'h0906: q0 = 16'hfff0; // 0x120c
	13'h0907: q0 = 16'h5240; // 0x120e
	13'h0908: q0 = 16'hd640; // 0x1210
	13'h0909: q0 = 16'h60d8; // 0x1212
	13'h090a: q0 = 16'h33c6; // 0x1214
	13'h090b: q0 = 16'h0001; // 0x1216
	13'h090c: q0 = 16'h893a; // 0x1218
	13'h090d: q0 = 16'h33c7; // 0x121a
	13'h090e: q0 = 16'h0001; // 0x121c
	13'h090f: q0 = 16'h7bd8; // 0x121e
	13'h0910: q0 = 16'hd779; // 0x1220
	13'h0911: q0 = 16'h0001; // 0x1222
	13'h0912: q0 = 16'h7594; // 0x1224
	13'h0913: q0 = 16'h0c79; // 0x1226
	13'h0914: q0 = 16'h0014; // 0x1228
	13'h0915: q0 = 16'h0001; // 0x122a
	13'h0916: q0 = 16'h7594; // 0x122c
	13'h0917: q0 = 16'h6f08; // 0x122e
	13'h0918: q0 = 16'h33fc; // 0x1230
	13'h0919: q0 = 16'h0014; // 0x1232
	13'h091a: q0 = 16'h0001; // 0x1234
	13'h091b: q0 = 16'h7594; // 0x1236
	13'h091c: q0 = 16'h3003; // 0x1238
	13'h091d: q0 = 16'h48c0; // 0x123a
	13'h091e: q0 = 16'hd1b9; // 0x123c
	13'h091f: q0 = 16'h0001; // 0x123e
	13'h0920: q0 = 16'h75aa; // 0x1240
	13'h0921: q0 = 16'h3003; // 0x1242
	13'h0922: q0 = 16'h48c0; // 0x1244
	13'h0923: q0 = 16'hd1b9; // 0x1246
	13'h0924: q0 = 16'h0001; // 0x1248
	13'h0925: q0 = 16'h75ce; // 0x124a
	13'h0926: q0 = 16'h4a43; // 0x124c
	13'h0927: q0 = 16'h670c; // 0x124e
	13'h0928: q0 = 16'h2ebc; // 0x1250
	13'h0929: q0 = 16'h0000; // 0x1252
	13'h092a: q0 = 16'hc53a; // 0x1254
	13'h092b: q0 = 16'h4eb9; // 0x1256
	13'h092c: q0 = 16'h0000; // 0x1258
	13'h092d: q0 = 16'h7e06; // 0x125a
	13'h092e: q0 = 16'h4a9f; // 0x125c
	13'h092f: q0 = 16'h4cdf; // 0x125e
	13'h0930: q0 = 16'h20f8; // 0x1260
	13'h0931: q0 = 16'h4e5e; // 0x1262
	13'h0932: q0 = 16'h4e75; // 0x1264
	13'h0933: q0 = 16'h4e56; // 0x1266
	13'h0934: q0 = 16'hfffc; // 0x1268
	13'h0935: q0 = 16'h4279; // 0x126a
	13'h0936: q0 = 16'h0001; // 0x126c
	13'h0937: q0 = 16'h7bd8; // 0x126e
	13'h0938: q0 = 16'h3039; // 0x1270
	13'h0939: q0 = 16'h0001; // 0x1272
	13'h093a: q0 = 16'h87dc; // 0x1274
	13'h093b: q0 = 16'h9179; // 0x1276
	13'h093c: q0 = 16'h0001; // 0x1278
	13'h093d: q0 = 16'h7594; // 0x127a
	13'h093e: q0 = 16'h4e5e; // 0x127c
	13'h093f: q0 = 16'h4e75; // 0x127e
	13'h0940: q0 = 16'h4e56; // 0x1280
	13'h0941: q0 = 16'h0000; // 0x1282
	13'h0942: q0 = 16'h48e7; // 0x1284
	13'h0943: q0 = 16'h1f00; // 0x1286
	13'h0944: q0 = 16'h3c2e; // 0x1288
	13'h0945: q0 = 16'h0008; // 0x128a
	13'h0946: q0 = 16'h3e2e; // 0x128c
	13'h0947: q0 = 16'h000a; // 0x128e
	13'h0948: q0 = 16'h3806; // 0x1290
	13'h0949: q0 = 16'hd87c; // 0x1292
	13'h094a: q0 = 16'h0012; // 0x1294
	13'h094b: q0 = 16'hb87c; // 0x1296
	13'h094c: q0 = 16'h0047; // 0x1298
	13'h094d: q0 = 16'h6f04; // 0x129a
	13'h094e: q0 = 16'h987c; // 0x129c
	13'h094f: q0 = 16'h0048; // 0x129e
	13'h0950: q0 = 16'h3e87; // 0x12a0
	13'h0951: q0 = 16'h3f04; // 0x12a2
	13'h0952: q0 = 16'h4eb9; // 0x12a4
	13'h0953: q0 = 16'h0000; // 0x12a6
	13'h0954: q0 = 16'ha730; // 0x12a8
	13'h0955: q0 = 16'h4a5f; // 0x12aa
	13'h0956: q0 = 16'h3a00; // 0x12ac
	13'h0957: q0 = 16'h3005; // 0x12ae
	13'h0958: q0 = 16'h4a9f; // 0x12b0
	13'h0959: q0 = 16'h4cdf; // 0x12b2
	13'h095a: q0 = 16'h00f0; // 0x12b4
	13'h095b: q0 = 16'h4e5e; // 0x12b6
	13'h095c: q0 = 16'h4e75; // 0x12b8
	13'h095d: q0 = 16'h4e56; // 0x12ba
	13'h095e: q0 = 16'hffdc; // 0x12bc
	13'h095f: q0 = 16'h48e7; // 0x12be
	13'h0960: q0 = 16'h1f04; // 0x12c0
	13'h0961: q0 = 16'h3839; // 0x12c2
	13'h0962: q0 = 16'h0001; // 0x12c4
	13'h0963: q0 = 16'h7594; // 0x12c6
	13'h0964: q0 = 16'h3c39; // 0x12c8
	13'h0965: q0 = 16'h0001; // 0x12ca
	13'h0966: q0 = 16'h758c; // 0x12cc
	13'h0967: q0 = 16'hb87c; // 0x12ce
	13'h0968: q0 = 16'h0001; // 0x12d0
	13'h0969: q0 = 16'h6f5e; // 0x12d2
	13'h096a: q0 = 16'h200e; // 0x12d4
	13'h096b: q0 = 16'hd0bc; // 0x12d6
	13'h096c: q0 = 16'hffff; // 0x12d8
	13'h096d: q0 = 16'hffe0; // 0x12da
	13'h096e: q0 = 16'h2e80; // 0x12dc
	13'h096f: q0 = 16'h3f04; // 0x12de
	13'h0970: q0 = 16'h4eb9; // 0x12e0
	13'h0971: q0 = 16'h0000; // 0x12e2
	13'h0972: q0 = 16'h0828; // 0x12e4
	13'h0973: q0 = 16'h4a5f; // 0x12e6
	13'h0974: q0 = 16'h2ebc; // 0x12e8
	13'h0975: q0 = 16'h0001; // 0x12ea
	13'h0976: q0 = 16'h8800; // 0x12ec
	13'h0977: q0 = 16'h200e; // 0x12ee
	13'h0978: q0 = 16'hd0bc; // 0x12f0
	13'h0979: q0 = 16'hffff; // 0x12f2
	13'h097a: q0 = 16'hffe0; // 0x12f4
	13'h097b: q0 = 16'h2f00; // 0x12f6
	13'h097c: q0 = 16'h4eb9; // 0x12f8
	13'h097d: q0 = 16'h0000; // 0x12fa
	13'h097e: q0 = 16'h0770; // 0x12fc
	13'h097f: q0 = 16'h4a9f; // 0x12fe
	13'h0980: q0 = 16'h41ee; // 0x1300
	13'h0981: q0 = 16'hffe0; // 0x1302
	13'h0982: q0 = 16'h23c8; // 0x1304
	13'h0983: q0 = 16'h0001; // 0x1306
	13'h0984: q0 = 16'h892a; // 0x1308
	13'h0985: q0 = 16'hbc7c; // 0x130a
	13'h0986: q0 = 16'h0001; // 0x130c
	13'h0987: q0 = 16'h6f16; // 0x130e
	13'h0988: q0 = 16'h23fc; // 0x1310
	13'h0989: q0 = 16'h0001; // 0x1312
	13'h098a: q0 = 16'h8840; // 0x1314
	13'h098b: q0 = 16'h0001; // 0x1316
	13'h098c: q0 = 16'h892e; // 0x1318
	13'h098d: q0 = 16'h23fc; // 0x131a
	13'h098e: q0 = 16'h0001; // 0x131c
	13'h098f: q0 = 16'h8820; // 0x131e
	13'h0990: q0 = 16'h0001; // 0x1320
	13'h0991: q0 = 16'h8932; // 0x1322
	13'h0992: q0 = 16'h600a; // 0x1324
	13'h0993: q0 = 16'h23fc; // 0x1326
	13'h0994: q0 = 16'h0001; // 0x1328
	13'h0995: q0 = 16'h8840; // 0x132a
	13'h0996: q0 = 16'h0001; // 0x132c
	13'h0997: q0 = 16'h8932; // 0x132e
	13'h0998: q0 = 16'h6026; // 0x1330
	13'h0999: q0 = 16'hb87c; // 0x1332
	13'h099a: q0 = 16'h0001; // 0x1334
	13'h099b: q0 = 16'h6616; // 0x1336
	13'h099c: q0 = 16'h23fc; // 0x1338
	13'h099d: q0 = 16'h0001; // 0x133a
	13'h099e: q0 = 16'h87e0; // 0x133c
	13'h099f: q0 = 16'h0001; // 0x133e
	13'h09a0: q0 = 16'h892a; // 0x1340
	13'h09a1: q0 = 16'h23fc; // 0x1342
	13'h09a2: q0 = 16'h0001; // 0x1344
	13'h09a3: q0 = 16'h8820; // 0x1346
	13'h09a4: q0 = 16'h0001; // 0x1348
	13'h09a5: q0 = 16'h8932; // 0x134a
	13'h09a6: q0 = 16'h600a; // 0x134c
	13'h09a7: q0 = 16'h23fc; // 0x134e
	13'h09a8: q0 = 16'h0001; // 0x1350
	13'h09a9: q0 = 16'h8860; // 0x1352
	13'h09aa: q0 = 16'h0001; // 0x1354
	13'h09ab: q0 = 16'h8932; // 0x1356
	13'h09ac: q0 = 16'h2d7c; // 0x1358
	13'h09ad: q0 = 16'h0000; // 0x135a
	13'h09ae: q0 = 16'h0008; // 0x135c
	13'h09af: q0 = 16'hffdc; // 0x135e
	13'h09b0: q0 = 16'h202e; // 0x1360
	13'h09b1: q0 = 16'hffdc; // 0x1362
	13'h09b2: q0 = 16'h4281; // 0x1364
	13'h09b3: q0 = 16'h7214; // 0x1366
	13'h09b4: q0 = 16'he3a0; // 0x1368
	13'h09b5: q0 = 16'h2d40; // 0x136a
	13'h09b6: q0 = 16'hffdc; // 0x136c
	13'h09b7: q0 = 16'h5cae; // 0x136e
	13'h09b8: q0 = 16'hffdc; // 0x1370
	13'h09b9: q0 = 16'h7e06; // 0x1372
	13'h09ba: q0 = 16'he947; // 0x1374
	13'h09bb: q0 = 16'hde7c; // 0x1376
	13'h09bc: q0 = 16'h000f; // 0x1378
	13'h09bd: q0 = 16'h3007; // 0x137a
	13'h09be: q0 = 16'he940; // 0x137c
	13'h09bf: q0 = 16'h48c0; // 0x137e
	13'h09c0: q0 = 16'hd1ae; // 0x1380
	13'h09c1: q0 = 16'hffdc; // 0x1382
	13'h09c2: q0 = 16'h202e; // 0x1384
	13'h09c3: q0 = 16'hffdc; // 0x1386
	13'h09c4: q0 = 16'h2040; // 0x1388
	13'h09c5: q0 = 16'h1e10; // 0x138a
	13'h09c6: q0 = 16'h4887; // 0x138c
	13'h09c7: q0 = 16'h52ae; // 0x138e
	13'h09c8: q0 = 16'hffdc; // 0x1390
	13'h09c9: q0 = 16'h202e; // 0x1392
	13'h09ca: q0 = 16'hffdc; // 0x1394
	13'h09cb: q0 = 16'h2040; // 0x1396
	13'h09cc: q0 = 16'h1010; // 0x1398
	13'h09cd: q0 = 16'h4880; // 0x139a
	13'h09ce: q0 = 16'h9047; // 0x139c
	13'h09cf: q0 = 16'hb07c; // 0x139e
	13'h09d0: q0 = 16'h002b; // 0x13a0
	13'h09d1: q0 = 16'h6708; // 0x13a2
	13'h09d2: q0 = 16'h33fc; // 0x13a4
	13'h09d3: q0 = 16'h0001; // 0x13a6
	13'h09d4: q0 = 16'h0001; // 0x13a8
	13'h09d5: q0 = 16'h7584; // 0x13aa
	13'h09d6: q0 = 16'h3a39; // 0x13ac
	13'h09d7: q0 = 16'h0001; // 0x13ae
	13'h09d8: q0 = 16'h893c; // 0x13b0
	13'h09d9: q0 = 16'h4247; // 0x13b2
	13'h09da: q0 = 16'h7c0f; // 0x13b4
	13'h09db: q0 = 16'h2a7c; // 0x13b6
	13'h09dc: q0 = 16'h0001; // 0x13b8
	13'h09dd: q0 = 16'h892a; // 0x13ba
	13'h09de: q0 = 16'hbe7c; // 0x13bc
	13'h09df: q0 = 16'h0003; // 0x13be
	13'h09e0: q0 = 16'h6c26; // 0x13c0
	13'h09e1: q0 = 16'hbc7c; // 0x13c2
	13'h09e2: q0 = 16'h0010; // 0x13c4
	13'h09e3: q0 = 16'h6602; // 0x13c6
	13'h09e4: q0 = 16'h5246; // 0x13c8
	13'h09e5: q0 = 16'h3e85; // 0x13ca
	13'h09e6: q0 = 16'h4267; // 0x13cc
	13'h09e7: q0 = 16'h3f3c; // 0x13ce
	13'h09e8: q0 = 16'h0064; // 0x13d0
	13'h09e9: q0 = 16'h3f06; // 0x13d2
	13'h09ea: q0 = 16'h2f15; // 0x13d4
	13'h09eb: q0 = 16'h4eb9; // 0x13d6
	13'h09ec: q0 = 16'h0000; // 0x13d8
	13'h09ed: q0 = 16'h026c; // 0x13da
	13'h09ee: q0 = 16'hdefc; // 0x13dc
	13'h09ef: q0 = 16'h000a; // 0x13de
	13'h09f0: q0 = 16'h5247; // 0x13e0
	13'h09f1: q0 = 16'h5246; // 0x13e2
	13'h09f2: q0 = 16'h588d; // 0x13e4
	13'h09f3: q0 = 16'h60d4; // 0x13e6
	13'h09f4: q0 = 16'h5245; // 0x13e8
	13'h09f5: q0 = 16'hba7c; // 0x13ea
	13'h09f6: q0 = 16'h003f; // 0x13ec
	13'h09f7: q0 = 16'h6f02; // 0x13ee
	13'h09f8: q0 = 16'h7a2d; // 0x13f0
	13'h09f9: q0 = 16'h33c5; // 0x13f2
	13'h09fa: q0 = 16'h0001; // 0x13f4
	13'h09fb: q0 = 16'h893c; // 0x13f6
	13'h09fc: q0 = 16'h4a9f; // 0x13f8
	13'h09fd: q0 = 16'h4cdf; // 0x13fa
	13'h09fe: q0 = 16'h20f0; // 0x13fc
	13'h09ff: q0 = 16'h4e5e; // 0x13fe
	13'h0a00: q0 = 16'h4e75; // 0x1400
	13'h0a01: q0 = 16'h4e56; // 0x1402
	13'h0a02: q0 = 16'hfffc; // 0x1404
	13'h0a03: q0 = 16'h48e7; // 0x1406
	13'h0a04: q0 = 16'h070c; // 0x1408
	13'h0a05: q0 = 16'h2a6e; // 0x140a
	13'h0a06: q0 = 16'h000a; // 0x140c
	13'h0a07: q0 = 16'h200e; // 0x140e
	13'h0a08: q0 = 16'hd0bc; // 0x1410
	13'h0a09: q0 = 16'hffff; // 0x1412
	13'h0a0a: q0 = 16'hfffc; // 0x1414
	13'h0a0b: q0 = 16'h2e80; // 0x1416
	13'h0a0c: q0 = 16'h3f2e; // 0x1418
	13'h0a0d: q0 = 16'h0008; // 0x141a
	13'h0a0e: q0 = 16'h4eb9; // 0x141c
	13'h0a0f: q0 = 16'h0000; // 0x141e
	13'h0a10: q0 = 16'h0828; // 0x1420
	13'h0a11: q0 = 16'h4a5f; // 0x1422
	13'h0a12: q0 = 16'h200e; // 0x1424
	13'h0a13: q0 = 16'hd0bc; // 0x1426
	13'h0a14: q0 = 16'hffff; // 0x1428
	13'h0a15: q0 = 16'hfffc; // 0x142a
	13'h0a16: q0 = 16'h2e80; // 0x142c
	13'h0a17: q0 = 16'h4eb9; // 0x142e
	13'h0a18: q0 = 16'h0000; // 0x1430
	13'h0a19: q0 = 16'h072e; // 0x1432
	13'h0a1a: q0 = 16'h3a80; // 0x1434
	13'h0a1b: q0 = 16'h302e; // 0x1436
	13'h0a1c: q0 = 16'h0012; // 0x1438
	13'h0a1d: q0 = 16'he740; // 0x143a
	13'h0a1e: q0 = 16'h48c0; // 0x143c
	13'h0a1f: q0 = 16'h2840; // 0x143e
	13'h0a20: q0 = 16'hd9fc; // 0x1440
	13'h0a21: q0 = 16'h0001; // 0x1442
	13'h0a22: q0 = 16'h75e8; // 0x1444
	13'h0a23: q0 = 16'h4247; // 0x1446
	13'h0a24: q0 = 16'hbe55; // 0x1448
	13'h0a25: q0 = 16'h6c48; // 0x144a
	13'h0a26: q0 = 16'h3207; // 0x144c
	13'h0a27: q0 = 16'h48c1; // 0x144e
	13'h0a28: q0 = 16'h200e; // 0x1450
	13'h0a29: q0 = 16'hd081; // 0x1452
	13'h0a2a: q0 = 16'h2040; // 0x1454
	13'h0a2b: q0 = 16'h1c28; // 0x1456
	13'h0a2c: q0 = 16'hfffc; // 0x1458
	13'h0a2d: q0 = 16'h4886; // 0x145a
	13'h0a2e: q0 = 16'hdc7c; // 0x145c
	13'h0a2f: q0 = 16'hffd0; // 0x145e
	13'h0a30: q0 = 16'h3006; // 0x1460
	13'h0a31: q0 = 16'h48c0; // 0x1462
	13'h0a32: q0 = 16'hd0bc; // 0x1464
	13'h0a33: q0 = 16'h0000; // 0x1466
	13'h0a34: q0 = 16'hc62e; // 0x1468
	13'h0a35: q0 = 16'h2040; // 0x146a
	13'h0a36: q0 = 16'h1c10; // 0x146c
	13'h0a37: q0 = 16'h4886; // 0x146e
	13'h0a38: q0 = 16'hcc7c; // 0x1470
	13'h0a39: q0 = 16'h00ff; // 0x1472
	13'h0a3a: q0 = 16'h3007; // 0x1474
	13'h0a3b: q0 = 16'he340; // 0x1476
	13'h0a3c: q0 = 16'h48c0; // 0x1478
	13'h0a3d: q0 = 16'hd08c; // 0x147a
	13'h0a3e: q0 = 16'h2040; // 0x147c
	13'h0a3f: q0 = 16'h3146; // 0x147e
	13'h0a40: q0 = 16'h0002; // 0x1480
	13'h0a41: q0 = 16'h3007; // 0x1482
	13'h0a42: q0 = 16'he340; // 0x1484
	13'h0a43: q0 = 16'h48c0; // 0x1486
	13'h0a44: q0 = 16'hd0ae; // 0x1488
	13'h0a45: q0 = 16'h000e; // 0x148a
	13'h0a46: q0 = 16'h2040; // 0x148c
	13'h0a47: q0 = 16'h3086; // 0x148e
	13'h0a48: q0 = 16'h5247; // 0x1490
	13'h0a49: q0 = 16'h60b4; // 0x1492
	13'h0a4a: q0 = 16'h0c55; // 0x1494
	13'h0a4b: q0 = 16'h0002; // 0x1496
	13'h0a4c: q0 = 16'h662c; // 0x1498
	13'h0a4d: q0 = 16'h206e; // 0x149a
	13'h0a4e: q0 = 16'h000e; // 0x149c
	13'h0a4f: q0 = 16'h3010; // 0x149e
	13'h0a50: q0 = 16'h226e; // 0x14a0
	13'h0a51: q0 = 16'h000e; // 0x14a2
	13'h0a52: q0 = 16'hb069; // 0x14a4
	13'h0a53: q0 = 16'h0002; // 0x14a6
	13'h0a54: q0 = 16'h6608; // 0x14a8
	13'h0a55: q0 = 16'h397c; // 0x14aa
	13'h0a56: q0 = 16'h0052; // 0x14ac
	13'h0a57: q0 = 16'h0006; // 0x14ae
	13'h0a58: q0 = 16'h600a; // 0x14b0
	13'h0a59: q0 = 16'h206e; // 0x14b2
	13'h0a5a: q0 = 16'h000e; // 0x14b4
	13'h0a5b: q0 = 16'h3968; // 0x14b6
	13'h0a5c: q0 = 16'h0002; // 0x14b8
	13'h0a5d: q0 = 16'h0006; // 0x14ba
	13'h0a5e: q0 = 16'h206e; // 0x14bc
	13'h0a5f: q0 = 16'h000e; // 0x14be
	13'h0a60: q0 = 16'h316c; // 0x14c0
	13'h0a61: q0 = 16'h0006; // 0x14c2
	13'h0a62: q0 = 16'h0004; // 0x14c4
	13'h0a63: q0 = 16'h4a9f; // 0x14c6
	13'h0a64: q0 = 16'h4cdf; // 0x14c8
	13'h0a65: q0 = 16'h30c0; // 0x14ca
	13'h0a66: q0 = 16'h4e5e; // 0x14cc
	13'h0a67: q0 = 16'h4e75; // 0x14ce
	13'h0a68: q0 = 16'h4e56; // 0x14d0
	13'h0a69: q0 = 16'hfffc; // 0x14d2
	13'h0a6a: q0 = 16'h48e7; // 0x14d4
	13'h0a6b: q0 = 16'h1f00; // 0x14d6
	13'h0a6c: q0 = 16'h3e2e; // 0x14d8
	13'h0a6d: q0 = 16'h0008; // 0x14da
	13'h0a6e: q0 = 16'h200e; // 0x14dc
	13'h0a6f: q0 = 16'hd0bc; // 0x14de
	13'h0a70: q0 = 16'hffff; // 0x14e0
	13'h0a71: q0 = 16'hfffc; // 0x14e2
	13'h0a72: q0 = 16'h2e80; // 0x14e4
	13'h0a73: q0 = 16'h3f07; // 0x14e6
	13'h0a74: q0 = 16'h4eb9; // 0x14e8
	13'h0a75: q0 = 16'h0000; // 0x14ea
	13'h0a76: q0 = 16'h0828; // 0x14ec
	13'h0a77: q0 = 16'h4a5f; // 0x14ee
	13'h0a78: q0 = 16'h4245; // 0x14f0
	13'h0a79: q0 = 16'h200e; // 0x14f2
	13'h0a7a: q0 = 16'hd0bc; // 0x14f4
	13'h0a7b: q0 = 16'hffff; // 0x14f6
	13'h0a7c: q0 = 16'hfffc; // 0x14f8
	13'h0a7d: q0 = 16'h2e80; // 0x14fa
	13'h0a7e: q0 = 16'h4eb9; // 0x14fc
	13'h0a7f: q0 = 16'h0000; // 0x14fe
	13'h0a80: q0 = 16'h072e; // 0x1500
	13'h0a81: q0 = 16'hb045; // 0x1502
	13'h0a82: q0 = 16'h6f54; // 0x1504
	13'h0a83: q0 = 16'h7c01; // 0x1506
	13'h0a84: q0 = 16'hbc7c; // 0x1508
	13'h0a85: q0 = 16'h0003; // 0x150a
	13'h0a86: q0 = 16'h6e48; // 0x150c
	13'h0a87: q0 = 16'h7003; // 0x150e
	13'h0a88: q0 = 16'h9046; // 0x1510
	13'h0a89: q0 = 16'hc1fc; // 0x1512
	13'h0a8a: q0 = 16'h000a; // 0x1514
	13'h0a8b: q0 = 16'h3800; // 0x1516
	13'h0a8c: q0 = 16'h3205; // 0x1518
	13'h0a8d: q0 = 16'h48c1; // 0x151a
	13'h0a8e: q0 = 16'h200e; // 0x151c
	13'h0a8f: q0 = 16'hd081; // 0x151e
	13'h0a90: q0 = 16'h2040; // 0x1520
	13'h0a91: q0 = 16'h1028; // 0x1522
	13'h0a92: q0 = 16'hfffc; // 0x1524
	13'h0a93: q0 = 16'h4880; // 0x1526
	13'h0a94: q0 = 16'hd07c; // 0x1528
	13'h0a95: q0 = 16'hffd0; // 0x152a
	13'h0a96: q0 = 16'hd840; // 0x152c
	13'h0a97: q0 = 16'h3005; // 0x152e
	13'h0a98: q0 = 16'he540; // 0x1530
	13'h0a99: q0 = 16'hd046; // 0x1532
	13'h0a9a: q0 = 16'he340; // 0x1534
	13'h0a9b: q0 = 16'h48c0; // 0x1536
	13'h0a9c: q0 = 16'hd0bc; // 0x1538
	13'h0a9d: q0 = 16'h0001; // 0x153a
	13'h0a9e: q0 = 16'h76f8; // 0x153c
	13'h0a9f: q0 = 16'h2040; // 0x153e
	13'h0aa0: q0 = 16'h3204; // 0x1540
	13'h0aa1: q0 = 16'h48c1; // 0x1542
	13'h0aa2: q0 = 16'hd2bc; // 0x1544
	13'h0aa3: q0 = 16'h0000; // 0x1546
	13'h0aa4: q0 = 16'hc62e; // 0x1548
	13'h0aa5: q0 = 16'h2241; // 0x154a
	13'h0aa6: q0 = 16'h1211; // 0x154c
	13'h0aa7: q0 = 16'h4881; // 0x154e
	13'h0aa8: q0 = 16'h3081; // 0x1550
	13'h0aa9: q0 = 16'h5246; // 0x1552
	13'h0aaa: q0 = 16'h60b2; // 0x1554
	13'h0aab: q0 = 16'h5245; // 0x1556
	13'h0aac: q0 = 16'h6098; // 0x1558
	13'h0aad: q0 = 16'h4a9f; // 0x155a
	13'h0aae: q0 = 16'h4cdf; // 0x155c
	13'h0aaf: q0 = 16'h00f0; // 0x155e
	13'h0ab0: q0 = 16'h4e5e; // 0x1560
	13'h0ab1: q0 = 16'h4e75; // 0x1562
	13'h0ab2: q0 = 16'h4e56; // 0x1564
	13'h0ab3: q0 = 16'h0000; // 0x1566
	13'h0ab4: q0 = 16'h48e7; // 0x1568
	13'h0ab5: q0 = 16'h0700; // 0x156a
	13'h0ab6: q0 = 16'h4247; // 0x156c
	13'h0ab7: q0 = 16'hbe7c; // 0x156e
	13'h0ab8: q0 = 16'h000a; // 0x1570
	13'h0ab9: q0 = 16'h6c00; // 0x1572
	13'h0aba: q0 = 16'h009c; // 0x1574
	13'h0abb: q0 = 16'h3007; // 0x1576
	13'h0abc: q0 = 16'h6000; // 0x1578
	13'h0abd: q0 = 16'h006c; // 0x157a
	13'h0abe: q0 = 16'h3c39; // 0x157c
	13'h0abf: q0 = 16'h0001; // 0x157e
	13'h0ac0: q0 = 16'h757a; // 0x1580
	13'h0ac1: q0 = 16'h5546; // 0x1582
	13'h0ac2: q0 = 16'h6000; // 0x1584
	13'h0ac3: q0 = 16'h0074; // 0x1586
	13'h0ac4: q0 = 16'h3c39; // 0x1588
	13'h0ac5: q0 = 16'h0001; // 0x158a
	13'h0ac6: q0 = 16'h757e; // 0x158c
	13'h0ac7: q0 = 16'h5346; // 0x158e
	13'h0ac8: q0 = 16'h6068; // 0x1590
	13'h0ac9: q0 = 16'h3039; // 0x1592
	13'h0aca: q0 = 16'h0001; // 0x1594
	13'h0acb: q0 = 16'h7580; // 0x1596
	13'h0acc: q0 = 16'h48c0; // 0x1598
	13'h0acd: q0 = 16'h81fc; // 0x159a
	13'h0ace: q0 = 16'h0032; // 0x159c
	13'h0acf: q0 = 16'h3c00; // 0x159e
	13'h0ad0: q0 = 16'h6058; // 0x15a0
	13'h0ad1: q0 = 16'h3039; // 0x15a2
	13'h0ad2: q0 = 16'h0001; // 0x15a4
	13'h0ad3: q0 = 16'h7582; // 0x15a6
	13'h0ad4: q0 = 16'h48c0; // 0x15a8
	13'h0ad5: q0 = 16'h81fc; // 0x15aa
	13'h0ad6: q0 = 16'h0032; // 0x15ac
	13'h0ad7: q0 = 16'h3c00; // 0x15ae
	13'h0ad8: q0 = 16'h6048; // 0x15b0
	13'h0ad9: q0 = 16'h3c39; // 0x15b2
	13'h0ada: q0 = 16'h0001; // 0x15b4
	13'h0adb: q0 = 16'h7586; // 0x15b6
	13'h0adc: q0 = 16'h6040; // 0x15b8
	13'h0add: q0 = 16'h3c39; // 0x15ba
	13'h0ade: q0 = 16'h0001; // 0x15bc
	13'h0adf: q0 = 16'h7588; // 0x15be
	13'h0ae0: q0 = 16'h6038; // 0x15c0
	13'h0ae1: q0 = 16'h3c39; // 0x15c2
	13'h0ae2: q0 = 16'h0001; // 0x15c4
	13'h0ae3: q0 = 16'h758a; // 0x15c6
	13'h0ae4: q0 = 16'h6030; // 0x15c8
	13'h0ae5: q0 = 16'h3c39; // 0x15ca
	13'h0ae6: q0 = 16'h0001; // 0x15cc
	13'h0ae7: q0 = 16'h758c; // 0x15ce
	13'h0ae8: q0 = 16'h6028; // 0x15d0
	13'h0ae9: q0 = 16'h3c39; // 0x15d2
	13'h0aea: q0 = 16'h0001; // 0x15d4
	13'h0aeb: q0 = 16'h758e; // 0x15d6
	13'h0aec: q0 = 16'h6020; // 0x15d8
	13'h0aed: q0 = 16'h3c39; // 0x15da
	13'h0aee: q0 = 16'h0001; // 0x15dc
	13'h0aef: q0 = 16'h7592; // 0x15de
	13'h0af0: q0 = 16'h5346; // 0x15e0
	13'h0af1: q0 = 16'h6016; // 0x15e2
	13'h0af2: q0 = 16'h6014; // 0x15e4
	13'h0af3: q0 = 16'hb07c; // 0x15e6
	13'h0af4: q0 = 16'h0009; // 0x15e8
	13'h0af5: q0 = 16'h620e; // 0x15ea
	13'h0af6: q0 = 16'he540; // 0x15ec
	13'h0af7: q0 = 16'h3040; // 0x15ee
	13'h0af8: q0 = 16'hd1fc; // 0x15f0
	13'h0af9: q0 = 16'h0000; // 0x15f2
	13'h0afa: q0 = 16'hc64c; // 0x15f4
	13'h0afb: q0 = 16'h2050; // 0x15f6
	13'h0afc: q0 = 16'h4ed0; // 0x15f8
	13'h0afd: q0 = 16'h3007; // 0x15fa
	13'h0afe: q0 = 16'he340; // 0x15fc
	13'h0aff: q0 = 16'h48c0; // 0x15fe
	13'h0b00: q0 = 16'hd0bc; // 0x1600
	13'h0b01: q0 = 16'h0001; // 0x1602
	13'h0b02: q0 = 16'h86b8; // 0x1604
	13'h0b03: q0 = 16'h2040; // 0x1606
	13'h0b04: q0 = 16'h3086; // 0x1608
	13'h0b05: q0 = 16'h5247; // 0x160a
	13'h0b06: q0 = 16'h6000; // 0x160c
	13'h0b07: q0 = 16'hff60; // 0x160e
	13'h0b08: q0 = 16'h4a9f; // 0x1610
	13'h0b09: q0 = 16'h4cdf; // 0x1612
	13'h0b0a: q0 = 16'h00c0; // 0x1614
	13'h0b0b: q0 = 16'h4e5e; // 0x1616
	13'h0b0c: q0 = 16'h4e75; // 0x1618
	13'h0b0d: q0 = 16'h4e56; // 0x161a
	13'h0b0e: q0 = 16'hfffc; // 0x161c
	13'h0b0f: q0 = 16'h48e7; // 0x161e
	13'h0b10: q0 = 16'h1f04; // 0x1620
	13'h0b11: q0 = 16'h2a6e; // 0x1622
	13'h0b12: q0 = 16'h0008; // 0x1624
	13'h0b13: q0 = 16'h3c3c; // 0x1626
	13'h0b14: q0 = 16'h0400; // 0x1628
	13'h0b15: q0 = 16'h4245; // 0x162a
	13'h0b16: q0 = 16'hba7c; // 0x162c
	13'h0b17: q0 = 16'h0004; // 0x162e
	13'h0b18: q0 = 16'h6c00; // 0x1630
	13'h0b19: q0 = 16'h0086; // 0x1632
	13'h0b1a: q0 = 16'h4a6d; // 0x1634
	13'h0b1b: q0 = 16'h0006; // 0x1636
	13'h0b1c: q0 = 16'h6f2c; // 0x1638
	13'h0b1d: q0 = 16'h302d; // 0x163a
	13'h0b1e: q0 = 16'h0004; // 0x163c
	13'h0b1f: q0 = 16'h5340; // 0x163e
	13'h0b20: q0 = 16'heb40; // 0x1640
	13'h0b21: q0 = 16'h322d; // 0x1642
	13'h0b22: q0 = 16'h0006; // 0x1644
	13'h0b23: q0 = 16'h5341; // 0x1646
	13'h0b24: q0 = 16'he541; // 0x1648
	13'h0b25: q0 = 16'hd041; // 0x164a
	13'h0b26: q0 = 16'h3e00; // 0x164c
	13'h0b27: q0 = 16'h3007; // 0x164e
	13'h0b28: q0 = 16'hd045; // 0x1650
	13'h0b29: q0 = 16'h48c0; // 0x1652
	13'h0b2a: q0 = 16'hd0bc; // 0x1654
	13'h0b2b: q0 = 16'h0000; // 0x1656
	13'h0b2c: q0 = 16'hf6ce; // 0x1658
	13'h0b2d: q0 = 16'h2040; // 0x165a
	13'h0b2e: q0 = 16'h1810; // 0x165c
	13'h0b2f: q0 = 16'h4884; // 0x165e
	13'h0b30: q0 = 16'hc87c; // 0x1660
	13'h0b31: q0 = 16'h00ff; // 0x1662
	13'h0b32: q0 = 16'h6002; // 0x1664
	13'h0b33: q0 = 16'h7840; // 0x1666
	13'h0b34: q0 = 16'h3d55; // 0x1668
	13'h0b35: q0 = 16'hfffe; // 0x166a
	13'h0b36: q0 = 16'h3d6d; // 0x166c
	13'h0b37: q0 = 16'h0002; // 0x166e
	13'h0b38: q0 = 16'hfffc; // 0x1670
	13'h0b39: q0 = 16'hba7c; // 0x1672
	13'h0b3a: q0 = 16'h0001; // 0x1674
	13'h0b3b: q0 = 16'h6706; // 0x1676
	13'h0b3c: q0 = 16'hba7c; // 0x1678
	13'h0b3d: q0 = 16'h0003; // 0x167a
	13'h0b3e: q0 = 16'h6604; // 0x167c
	13'h0b3f: q0 = 16'hdd6e; // 0x167e
	13'h0b40: q0 = 16'hfffe; // 0x1680
	13'h0b41: q0 = 16'hba7c; // 0x1682
	13'h0b42: q0 = 16'h0002; // 0x1684
	13'h0b43: q0 = 16'h6c04; // 0x1686
	13'h0b44: q0 = 16'hdd6e; // 0x1688
	13'h0b45: q0 = 16'hfffc; // 0x168a
	13'h0b46: q0 = 16'h302d; // 0x168c
	13'h0b47: q0 = 16'h0004; // 0x168e
	13'h0b48: q0 = 16'h5340; // 0x1690
	13'h0b49: q0 = 16'he340; // 0x1692
	13'h0b4a: q0 = 16'h48c0; // 0x1694
	13'h0b4b: q0 = 16'hd0bc; // 0x1696
	13'h0b4c: q0 = 16'h0000; // 0x1698
	13'h0b4d: q0 = 16'hf6c4; // 0x169a
	13'h0b4e: q0 = 16'h2040; // 0x169c
	13'h0b4f: q0 = 16'h3e90; // 0x169e
	13'h0b50: q0 = 16'h3f04; // 0x16a0
	13'h0b51: q0 = 16'h3f2e; // 0x16a2
	13'h0b52: q0 = 16'hfffc; // 0x16a4
	13'h0b53: q0 = 16'h3f2e; // 0x16a6
	13'h0b54: q0 = 16'hfffe; // 0x16a8
	13'h0b55: q0 = 16'h4eb9; // 0x16aa
	13'h0b56: q0 = 16'h0000; // 0x16ac
	13'h0b57: q0 = 16'h3f80; // 0x16ae
	13'h0b58: q0 = 16'h5c4f; // 0x16b0
	13'h0b59: q0 = 16'h5245; // 0x16b2
	13'h0b5a: q0 = 16'h6000; // 0x16b4
	13'h0b5b: q0 = 16'hff76; // 0x16b6
	13'h0b5c: q0 = 16'h4a9f; // 0x16b8
	13'h0b5d: q0 = 16'h4cdf; // 0x16ba
	13'h0b5e: q0 = 16'h20f0; // 0x16bc
	13'h0b5f: q0 = 16'h4e5e; // 0x16be
	13'h0b60: q0 = 16'h4e75; // 0x16c0
	13'h0b61: q0 = 16'h4e56; // 0x16c2
	13'h0b62: q0 = 16'h0000; // 0x16c4
	13'h0b63: q0 = 16'h48e7; // 0x16c6
	13'h0b64: q0 = 16'h0304; // 0x16c8
	13'h0b65: q0 = 16'h2a7c; // 0x16ca
	13'h0b66: q0 = 16'h0001; // 0x16cc
	13'h0b67: q0 = 16'h89be; // 0x16ce
	13'h0b68: q0 = 16'h4247; // 0x16d0
	13'h0b69: q0 = 16'hbe79; // 0x16d2
	13'h0b6a: q0 = 16'h0001; // 0x16d4
	13'h0b6b: q0 = 16'h7fbc; // 0x16d6
	13'h0b6c: q0 = 16'h6c2a; // 0x16d8
	13'h0b6d: q0 = 16'h302d; // 0x16da
	13'h0b6e: q0 = 16'h000e; // 0x16dc
	13'h0b6f: q0 = 16'hc07c; // 0x16de
	13'h0b70: q0 = 16'h000f; // 0x16e0
	13'h0b71: q0 = 16'hb07c; // 0x16e2
	13'h0b72: q0 = 16'h0003; // 0x16e4
	13'h0b73: q0 = 16'h670e; // 0x16e6
	13'h0b74: q0 = 16'h302d; // 0x16e8
	13'h0b75: q0 = 16'h000e; // 0x16ea
	13'h0b76: q0 = 16'hc07c; // 0x16ec
	13'h0b77: q0 = 16'h000f; // 0x16ee
	13'h0b78: q0 = 16'hb07c; // 0x16f0
	13'h0b79: q0 = 16'h0004; // 0x16f2
	13'h0b7a: q0 = 16'h6604; // 0x16f4
	13'h0b7b: q0 = 16'h4240; // 0x16f6
	13'h0b7c: q0 = 16'h600c; // 0x16f8
	13'h0b7d: q0 = 16'hdbfc; // 0x16fa
	13'h0b7e: q0 = 16'h0000; // 0x16fc
	13'h0b7f: q0 = 16'h002e; // 0x16fe
	13'h0b80: q0 = 16'h5247; // 0x1700
	13'h0b81: q0 = 16'h60ce; // 0x1702
	13'h0b82: q0 = 16'h7001; // 0x1704
	13'h0b83: q0 = 16'h4a9f; // 0x1706
	13'h0b84: q0 = 16'h4cdf; // 0x1708
	13'h0b85: q0 = 16'h2080; // 0x170a
	13'h0b86: q0 = 16'h4e5e; // 0x170c
	13'h0b87: q0 = 16'h4e75; // 0x170e
	13'h0b88: q0 = 16'h4e56; // 0x1710
	13'h0b89: q0 = 16'h0000; // 0x1712
	13'h0b8a: q0 = 16'h48e7; // 0x1714
	13'h0b8b: q0 = 16'h0304; // 0x1716
	13'h0b8c: q0 = 16'h4a6e; // 0x1718
	13'h0b8d: q0 = 16'h0008; // 0x171a
	13'h0b8e: q0 = 16'h6600; // 0x171c
	13'h0b8f: q0 = 16'h008a; // 0x171e
	13'h0b90: q0 = 16'h4eb9; // 0x1720
	13'h0b91: q0 = 16'h0000; // 0x1722
	13'h0b92: q0 = 16'h1e8a; // 0x1724
	13'h0b93: q0 = 16'h33fc; // 0x1726
	13'h0b94: q0 = 16'h0004; // 0x1728
	13'h0b95: q0 = 16'h0001; // 0x172a
	13'h0b96: q0 = 16'h7fbc; // 0x172c
	13'h0b97: q0 = 16'h2a7c; // 0x172e
	13'h0b98: q0 = 16'h0001; // 0x1730
	13'h0b99: q0 = 16'h89be; // 0x1732
	13'h0b9a: q0 = 16'h4247; // 0x1734
	13'h0b9b: q0 = 16'hbe79; // 0x1736
	13'h0b9c: q0 = 16'h0001; // 0x1738
	13'h0b9d: q0 = 16'h7fbc; // 0x173a
	13'h0b9e: q0 = 16'h6c66; // 0x173c
	13'h0b9f: q0 = 16'h426d; // 0x173e
	13'h0ba0: q0 = 16'h000e; // 0x1740
	13'h0ba1: q0 = 16'h302d; // 0x1742
	13'h0ba2: q0 = 16'h000e; // 0x1744
	13'h0ba3: q0 = 16'hc07c; // 0x1746
	13'h0ba4: q0 = 16'hf0f0; // 0x1748
	13'h0ba5: q0 = 16'h807c; // 0x174a
	13'h0ba6: q0 = 16'h0002; // 0x174c
	13'h0ba7: q0 = 16'h3b40; // 0x174e
	13'h0ba8: q0 = 16'h000e; // 0x1750
	13'h0ba9: q0 = 16'h2b7c; // 0x1752
	13'h0baa: q0 = 16'h0000; // 0x1754
	13'h0bab: q0 = 16'h2710; // 0x1756
	13'h0bac: q0 = 16'h002a; // 0x1758
	13'h0bad: q0 = 16'h4255; // 0x175a
	13'h0bae: q0 = 16'h42ad; // 0x175c
	13'h0baf: q0 = 16'h0010; // 0x175e
	13'h0bb0: q0 = 16'h3007; // 0x1760
	13'h0bb1: q0 = 16'hc1fc; // 0x1762
	13'h0bb2: q0 = 16'h0006; // 0x1764
	13'h0bb3: q0 = 16'hd0bc; // 0x1766
	13'h0bb4: q0 = 16'h0000; // 0x1768
	13'h0bb5: q0 = 16'hc868; // 0x176a
	13'h0bb6: q0 = 16'h2b40; // 0x176c
	13'h0bb7: q0 = 16'h001a; // 0x176e
	13'h0bb8: q0 = 16'h206d; // 0x1770
	13'h0bb9: q0 = 16'h001a; // 0x1772
	13'h0bba: q0 = 16'h3010; // 0x1774
	13'h0bbb: q0 = 16'h5340; // 0x1776
	13'h0bbc: q0 = 16'hc1fc; // 0x1778
	13'h0bbd: q0 = 16'h000b; // 0x177a
	13'h0bbe: q0 = 16'h48c0; // 0x177c
	13'h0bbf: q0 = 16'hd0bc; // 0x177e
	13'h0bc0: q0 = 16'h0000; // 0x1780
	13'h0bc1: q0 = 16'hc89c; // 0x1782
	13'h0bc2: q0 = 16'h226d; // 0x1784
	13'h0bc3: q0 = 16'h001a; // 0x1786
	13'h0bc4: q0 = 16'h3211; // 0x1788
	13'h0bc5: q0 = 16'h5341; // 0x178a
	13'h0bc6: q0 = 16'he541; // 0x178c
	13'h0bc7: q0 = 16'h48c1; // 0x178e
	13'h0bc8: q0 = 16'hd2bc; // 0x1790
	13'h0bc9: q0 = 16'h0001; // 0x1792
	13'h0bca: q0 = 16'h85fe; // 0x1794
	13'h0bcb: q0 = 16'h2241; // 0x1796
	13'h0bcc: q0 = 16'h2280; // 0x1798
	13'h0bcd: q0 = 16'hdbfc; // 0x179a
	13'h0bce: q0 = 16'h0000; // 0x179c
	13'h0bcf: q0 = 16'h002e; // 0x179e
	13'h0bd0: q0 = 16'h5247; // 0x17a0
	13'h0bd1: q0 = 16'h6092; // 0x17a2
	13'h0bd2: q0 = 16'h6000; // 0x17a4
	13'h0bd3: q0 = 16'h007a; // 0x17a6
	13'h0bd4: q0 = 16'h0c6e; // 0x17a8
	13'h0bd5: q0 = 16'h0002; // 0x17aa
	13'h0bd6: q0 = 16'h0008; // 0x17ac
	13'h0bd7: q0 = 16'h6628; // 0x17ae
	13'h0bd8: q0 = 16'h2a7c; // 0x17b0
	13'h0bd9: q0 = 16'h0001; // 0x17b2
	13'h0bda: q0 = 16'h89be; // 0x17b4
	13'h0bdb: q0 = 16'h4247; // 0x17b6
	13'h0bdc: q0 = 16'hbe79; // 0x17b8
	13'h0bdd: q0 = 16'h0001; // 0x17ba
	13'h0bde: q0 = 16'h7fbc; // 0x17bc
	13'h0bdf: q0 = 16'h6c16; // 0x17be
	13'h0be0: q0 = 16'h426d; // 0x17c0
	13'h0be1: q0 = 16'h000e; // 0x17c2
	13'h0be2: q0 = 16'h2e8d; // 0x17c4
	13'h0be3: q0 = 16'h4eb9; // 0x17c6
	13'h0be4: q0 = 16'h0000; // 0x17c8
	13'h0be5: q0 = 16'h1f50; // 0x17ca
	13'h0be6: q0 = 16'hdbfc; // 0x17cc
	13'h0be7: q0 = 16'h0000; // 0x17ce
	13'h0be8: q0 = 16'h002e; // 0x17d0
	13'h0be9: q0 = 16'h5247; // 0x17d2
	13'h0bea: q0 = 16'h60e2; // 0x17d4
	13'h0beb: q0 = 16'h6048; // 0x17d6
	13'h0bec: q0 = 16'h0c6e; // 0x17d8
	13'h0bed: q0 = 16'h0005; // 0x17da
	13'h0bee: q0 = 16'h0008; // 0x17dc
	13'h0bef: q0 = 16'h6640; // 0x17de
	13'h0bf0: q0 = 16'h2a7c; // 0x17e0
	13'h0bf1: q0 = 16'h0001; // 0x17e2
	13'h0bf2: q0 = 16'h89be; // 0x17e4
	13'h0bf3: q0 = 16'h4247; // 0x17e6
	13'h0bf4: q0 = 16'hbe79; // 0x17e8
	13'h0bf5: q0 = 16'h0001; // 0x17ea
	13'h0bf6: q0 = 16'h7fbc; // 0x17ec
	13'h0bf7: q0 = 16'h6c1c; // 0x17ee
	13'h0bf8: q0 = 16'h42ad; // 0x17f0
	13'h0bf9: q0 = 16'h002a; // 0x17f2
	13'h0bfa: q0 = 16'h3e87; // 0x17f4
	13'h0bfb: q0 = 16'h5257; // 0x17f6
	13'h0bfc: q0 = 16'h2f0d; // 0x17f8
	13'h0bfd: q0 = 16'h4eb9; // 0x17fa
	13'h0bfe: q0 = 16'h0000; // 0x17fc
	13'h0bff: q0 = 16'h2c02; // 0x17fe
	13'h0c00: q0 = 16'h4a9f; // 0x1800
	13'h0c01: q0 = 16'hdbfc; // 0x1802
	13'h0c02: q0 = 16'h0000; // 0x1804
	13'h0c03: q0 = 16'h002e; // 0x1806
	13'h0c04: q0 = 16'h5247; // 0x1808
	13'h0c05: q0 = 16'h60dc; // 0x180a
	13'h0c06: q0 = 16'h7041; // 0x180c
	13'h0c07: q0 = 16'h2279; // 0x180e
	13'h0c08: q0 = 16'h0001; // 0x1810
	13'h0c09: q0 = 16'h7fb8; // 0x1812
	13'h0c0a: q0 = 16'h3211; // 0x1814
	13'h0c0b: q0 = 16'he541; // 0x1816
	13'h0c0c: q0 = 16'h9041; // 0x1818
	13'h0c0d: q0 = 16'h33c0; // 0x181a
	13'h0c0e: q0 = 16'h0001; // 0x181c
	13'h0c0f: q0 = 16'h7f28; // 0x181e
	13'h0c10: q0 = 16'h4a9f; // 0x1820
	13'h0c11: q0 = 16'h4cdf; // 0x1822
	13'h0c12: q0 = 16'h2080; // 0x1824
	13'h0c13: q0 = 16'h4e5e; // 0x1826
	13'h0c14: q0 = 16'h4e75; // 0x1828
	13'h0c15: q0 = 16'h4e56; // 0x182a
	13'h0c16: q0 = 16'hfffa; // 0x182c
	13'h0c17: q0 = 16'h48e7; // 0x182e
	13'h0c18: q0 = 16'h0104; // 0x1830
	13'h0c19: q0 = 16'h2a7c; // 0x1832
	13'h0c1a: q0 = 16'h0001; // 0x1834
	13'h0c1b: q0 = 16'h89be; // 0x1836
	13'h0c1c: q0 = 16'h426e; // 0x1838
	13'h0c1d: q0 = 16'hfffe; // 0x183a
	13'h0c1e: q0 = 16'h302e; // 0x183c
	13'h0c1f: q0 = 16'hfffe; // 0x183e
	13'h0c20: q0 = 16'hb079; // 0x1840
	13'h0c21: q0 = 16'h0001; // 0x1842
	13'h0c22: q0 = 16'h7fbc; // 0x1844
	13'h0c23: q0 = 16'h6c30; // 0x1846
	13'h0c24: q0 = 16'h302d; // 0x1848
	13'h0c25: q0 = 16'h000e; // 0x184a
	13'h0c26: q0 = 16'hc07c; // 0x184c
	13'h0c27: q0 = 16'h000f; // 0x184e
	13'h0c28: q0 = 16'h661a; // 0x1850
	13'h0c29: q0 = 16'h206e; // 0x1852
	13'h0c2a: q0 = 16'h0008; // 0x1854
	13'h0c2b: q0 = 16'h226d; // 0x1856
	13'h0c2c: q0 = 16'h001e; // 0x1858
	13'h0c2d: q0 = 16'h3091; // 0x185a
	13'h0c2e: q0 = 16'h206e; // 0x185c
	13'h0c2f: q0 = 16'h000c; // 0x185e
	13'h0c30: q0 = 16'h226d; // 0x1860
	13'h0c31: q0 = 16'h001e; // 0x1862
	13'h0c32: q0 = 16'h30a9; // 0x1864
	13'h0c33: q0 = 16'h0002; // 0x1866
	13'h0c34: q0 = 16'h7001; // 0x1868
	13'h0c35: q0 = 16'h605a; // 0x186a
	13'h0c36: q0 = 16'hdbfc; // 0x186c
	13'h0c37: q0 = 16'h0000; // 0x186e
	13'h0c38: q0 = 16'h002e; // 0x1870
	13'h0c39: q0 = 16'h526e; // 0x1872
	13'h0c3a: q0 = 16'hfffe; // 0x1874
	13'h0c3b: q0 = 16'h60c4; // 0x1876
	13'h0c3c: q0 = 16'h2d7c; // 0x1878
	13'h0c3d: q0 = 16'h0000; // 0x187a
	13'h0c3e: q0 = 16'h0001; // 0x187c
	13'h0c3f: q0 = 16'hfffa; // 0x187e
	13'h0c40: q0 = 16'h202e; // 0x1880
	13'h0c41: q0 = 16'hfffa; // 0x1882
	13'h0c42: q0 = 16'h4281; // 0x1884
	13'h0c43: q0 = 16'h7217; // 0x1886
	13'h0c44: q0 = 16'he3a0; // 0x1888
	13'h0c45: q0 = 16'h2d40; // 0x188a
	13'h0c46: q0 = 16'hfffa; // 0x188c
	13'h0c47: q0 = 16'h06ae; // 0x188e
	13'h0c48: q0 = 16'h0000; // 0x1890
	13'h0c49: q0 = 16'h0706; // 0x1892
	13'h0c4a: q0 = 16'hfffa; // 0x1894
	13'h0c4b: q0 = 16'h06ae; // 0x1896
	13'h0c4c: q0 = 16'h0000; // 0x1898
	13'h0c4d: q0 = 16'h0030; // 0x189a
	13'h0c4e: q0 = 16'hfffa; // 0x189c
	13'h0c4f: q0 = 16'h202e; // 0x189e
	13'h0c50: q0 = 16'hfffa; // 0x18a0
	13'h0c51: q0 = 16'h2040; // 0x18a2
	13'h0c52: q0 = 16'h1028; // 0x18a4
	13'h0c53: q0 = 16'h0001; // 0x18a6
	13'h0c54: q0 = 16'h4880; // 0x18a8
	13'h0c55: q0 = 16'h222e; // 0x18aa
	13'h0c56: q0 = 16'hfffa; // 0x18ac
	13'h0c57: q0 = 16'h2241; // 0x18ae
	13'h0c58: q0 = 16'h1211; // 0x18b0
	13'h0c59: q0 = 16'h4881; // 0x18b2
	13'h0c5a: q0 = 16'hd041; // 0x18b4
	13'h0c5b: q0 = 16'hb07c; // 0x18b6
	13'h0c5c: q0 = 16'h006a; // 0x18b8
	13'h0c5d: q0 = 16'h6708; // 0x18ba
	13'h0c5e: q0 = 16'h33fc; // 0x18bc
	13'h0c5f: q0 = 16'h0001; // 0x18be
	13'h0c60: q0 = 16'h0001; // 0x18c0
	13'h0c61: q0 = 16'h7590; // 0x18c2
	13'h0c62: q0 = 16'h4240; // 0x18c4
	13'h0c63: q0 = 16'h4a9f; // 0x18c6
	13'h0c64: q0 = 16'h4cdf; // 0x18c8
	13'h0c65: q0 = 16'h2000; // 0x18ca
	13'h0c66: q0 = 16'h4e5e; // 0x18cc
	13'h0c67: q0 = 16'h4e75; // 0x18ce
	13'h0c68: q0 = 16'h4e56; // 0x18d0
	13'h0c69: q0 = 16'hfffc; // 0x18d2
	13'h0c6a: q0 = 16'h48e7; // 0x18d4
	13'h0c6b: q0 = 16'h0f04; // 0x18d6
	13'h0c6c: q0 = 16'h2a7c; // 0x18d8
	13'h0c6d: q0 = 16'h0001; // 0x18da
	13'h0c6e: q0 = 16'h89be; // 0x18dc
	13'h0c6f: q0 = 16'h4247; // 0x18de
	13'h0c70: q0 = 16'hbe79; // 0x18e0
	13'h0c71: q0 = 16'h0001; // 0x18e2
	13'h0c72: q0 = 16'h7fbc; // 0x18e4
	13'h0c73: q0 = 16'h6c14; // 0x18e6
	13'h0c74: q0 = 16'h4aad; // 0x18e8
	13'h0c75: q0 = 16'h002a; // 0x18ea
	13'h0c76: q0 = 16'h6f04; // 0x18ec
	13'h0c77: q0 = 16'h53ad; // 0x18ee
	13'h0c78: q0 = 16'h002a; // 0x18f0
	13'h0c79: q0 = 16'hdbfc; // 0x18f2
	13'h0c7a: q0 = 16'h0000; // 0x18f4
	13'h0c7b: q0 = 16'h002e; // 0x18f6
	13'h0c7c: q0 = 16'h5247; // 0x18f8
	13'h0c7d: q0 = 16'h60e4; // 0x18fa
	13'h0c7e: q0 = 16'h2a7c; // 0x18fc
	13'h0c7f: q0 = 16'h0001; // 0x18fe
	13'h0c80: q0 = 16'h89be; // 0x1900
	13'h0c81: q0 = 16'h4247; // 0x1902
	13'h0c82: q0 = 16'hbe79; // 0x1904
	13'h0c83: q0 = 16'h0001; // 0x1906
	13'h0c84: q0 = 16'h7fbc; // 0x1908
	13'h0c85: q0 = 16'h6c00; // 0x190a
	13'h0c86: q0 = 16'h04ee; // 0x190c
	13'h0c87: q0 = 16'h302d; // 0x190e
	13'h0c88: q0 = 16'h000e; // 0x1910
	13'h0c89: q0 = 16'hc07c; // 0x1912
	13'h0c8a: q0 = 16'h000f; // 0x1914
	13'h0c8b: q0 = 16'hb07c; // 0x1916
	13'h0c8c: q0 = 16'h0002; // 0x1918
	13'h0c8d: q0 = 16'h671c; // 0x191a
	13'h0c8e: q0 = 16'h302d; // 0x191c
	13'h0c8f: q0 = 16'h000e; // 0x191e
	13'h0c90: q0 = 16'hc07c; // 0x1920
	13'h0c91: q0 = 16'h000f; // 0x1922
	13'h0c92: q0 = 16'hb07c; // 0x1924
	13'h0c93: q0 = 16'h0003; // 0x1926
	13'h0c94: q0 = 16'h670e; // 0x1928
	13'h0c95: q0 = 16'h302d; // 0x192a
	13'h0c96: q0 = 16'h000e; // 0x192c
	13'h0c97: q0 = 16'hc07c; // 0x192e
	13'h0c98: q0 = 16'h000f; // 0x1930
	13'h0c99: q0 = 16'hb07c; // 0x1932
	13'h0c9a: q0 = 16'h0004; // 0x1934
	13'h0c9b: q0 = 16'h660c; // 0x1936
	13'h0c9c: q0 = 16'h2e8d; // 0x1938
	13'h0c9d: q0 = 16'h4eb9; // 0x193a
	13'h0c9e: q0 = 16'h0000; // 0x193c
	13'h0c9f: q0 = 16'h291a; // 0x193e
	13'h0ca0: q0 = 16'h6000; // 0x1940
	13'h0ca1: q0 = 16'h04ac; // 0x1942
	13'h0ca2: q0 = 16'h4eb9; // 0x1944
	13'h0ca3: q0 = 16'h0000; // 0x1946
	13'h0ca4: q0 = 16'h4738; // 0x1948
	13'h0ca5: q0 = 16'hb07c; // 0x194a
	13'h0ca6: q0 = 16'h0002; // 0x194c
	13'h0ca7: q0 = 16'h662a; // 0x194e
	13'h0ca8: q0 = 16'h206d; // 0x1950
	13'h0ca9: q0 = 16'h001e; // 0x1952
	13'h0caa: q0 = 16'h317c; // 0x1954
	13'h0cab: q0 = 16'h0017; // 0x1956
	13'h0cac: q0 = 16'h0006; // 0x1958
	13'h0cad: q0 = 16'h3e95; // 0x195a
	13'h0cae: q0 = 16'h202d; // 0x195c
	13'h0caf: q0 = 16'h001e; // 0x195e
	13'h0cb0: q0 = 16'h5c80; // 0x1960
	13'h0cb1: q0 = 16'h2f00; // 0x1962
	13'h0cb2: q0 = 16'h4eb9; // 0x1964
	13'h0cb3: q0 = 16'h0000; // 0x1966
	13'h0cb4: q0 = 16'h3ee6; // 0x1968
	13'h0cb5: q0 = 16'h4a9f; // 0x196a
	13'h0cb6: q0 = 16'h206d; // 0x196c
	13'h0cb7: q0 = 16'h0026; // 0x196e
	13'h0cb8: q0 = 16'h317c; // 0x1970
	13'h0cb9: q0 = 16'h0017; // 0x1972
	13'h0cba: q0 = 16'h0006; // 0x1974
	13'h0cbb: q0 = 16'h6000; // 0x1976
	13'h0cbc: q0 = 16'h0476; // 0x1978
	13'h0cbd: q0 = 16'h4eb9; // 0x197a
	13'h0cbe: q0 = 16'h0000; // 0x197c
	13'h0cbf: q0 = 16'h4ec6; // 0x197e
	13'h0cc0: q0 = 16'hb07c; // 0x1980
	13'h0cc1: q0 = 16'h0006; // 0x1982
	13'h0cc2: q0 = 16'h6716; // 0x1984
	13'h0cc3: q0 = 16'h4eb9; // 0x1986
	13'h0cc4: q0 = 16'h0000; // 0x1988
	13'h0cc5: q0 = 16'h4ec6; // 0x198a
	13'h0cc6: q0 = 16'h4a40; // 0x198c
	13'h0cc7: q0 = 16'h6f58; // 0x198e
	13'h0cc8: q0 = 16'h4eb9; // 0x1990
	13'h0cc9: q0 = 16'h0000; // 0x1992
	13'h0cca: q0 = 16'h4ec6; // 0x1994
	13'h0ccb: q0 = 16'hb07c; // 0x1996
	13'h0ccc: q0 = 16'h0005; // 0x1998
	13'h0ccd: q0 = 16'h6c4c; // 0x199a
	13'h0cce: q0 = 16'h082d; // 0x199c
	13'h0ccf: q0 = 16'h0004; // 0x199e
	13'h0cd0: q0 = 16'h000f; // 0x19a0
	13'h0cd1: q0 = 16'h6644; // 0x19a2
	13'h0cd2: q0 = 16'h3b7c; // 0x19a4
	13'h0cd3: q0 = 16'h0001; // 0x19a6
	13'h0cd4: q0 = 16'h000c; // 0x19a8
	13'h0cd5: q0 = 16'h426d; // 0x19aa
	13'h0cd6: q0 = 16'h000a; // 0x19ac
	13'h0cd7: q0 = 16'h082d; // 0x19ae
	13'h0cd8: q0 = 16'h0000; // 0x19b0
	13'h0cd9: q0 = 16'h000e; // 0x19b2
	13'h0cda: q0 = 16'h670c; // 0x19b4
	13'h0cdb: q0 = 16'h302d; // 0x19b6
	13'h0cdc: q0 = 16'h000e; // 0x19b8
	13'h0cdd: q0 = 16'hc07c; // 0x19ba
	13'h0cde: q0 = 16'hfeff; // 0x19bc
	13'h0cdf: q0 = 16'h3b40; // 0x19be
	13'h0ce0: q0 = 16'h000e; // 0x19c0
	13'h0ce1: q0 = 16'h082d; // 0x19c2
	13'h0ce2: q0 = 16'h0001; // 0x19c4
	13'h0ce3: q0 = 16'h000e; // 0x19c6
	13'h0ce4: q0 = 16'h670c; // 0x19c8
	13'h0ce5: q0 = 16'h302d; // 0x19ca
	13'h0ce6: q0 = 16'h000e; // 0x19cc
	13'h0ce7: q0 = 16'hc07c; // 0x19ce
	13'h0ce8: q0 = 16'hfdff; // 0x19d0
	13'h0ce9: q0 = 16'h3b40; // 0x19d2
	13'h0cea: q0 = 16'h000e; // 0x19d4
	13'h0ceb: q0 = 16'h426d; // 0x19d6
	13'h0cec: q0 = 16'h0002; // 0x19d8
	13'h0ced: q0 = 16'h426d; // 0x19da
	13'h0cee: q0 = 16'h0004; // 0x19dc
	13'h0cef: q0 = 16'h426d; // 0x19de
	13'h0cf0: q0 = 16'h0006; // 0x19e0
	13'h0cf1: q0 = 16'h006d; // 0x19e2
	13'h0cf2: q0 = 16'h0010; // 0x19e4
	13'h0cf3: q0 = 16'h000e; // 0x19e6
	13'h0cf4: q0 = 16'h4a79; // 0x19e8
	13'h0cf5: q0 = 16'h0001; // 0x19ea
	13'h0cf6: q0 = 16'h7f2a; // 0x19ec
	13'h0cf7: q0 = 16'h6642; // 0x19ee
	13'h0cf8: q0 = 16'h302d; // 0x19f0
	13'h0cf9: q0 = 16'h000e; // 0x19f2
	13'h0cfa: q0 = 16'hc07c; // 0x19f4
	13'h0cfb: q0 = 16'h000f; // 0x19f6
	13'h0cfc: q0 = 16'h670e; // 0x19f8
	13'h0cfd: q0 = 16'h302d; // 0x19fa
	13'h0cfe: q0 = 16'h000e; // 0x19fc
	13'h0cff: q0 = 16'hc07c; // 0x19fe
	13'h0d00: q0 = 16'h000f; // 0x1a00
	13'h0d01: q0 = 16'hb07c; // 0x1a02
	13'h0d02: q0 = 16'h0001; // 0x1a04
	13'h0d03: q0 = 16'h662a; // 0x1a06
	13'h0d04: q0 = 16'h2e8d; // 0x1a08
	13'h0d05: q0 = 16'h4eb9; // 0x1a0a
	13'h0d06: q0 = 16'h0000; // 0x1a0c
	13'h0d07: q0 = 16'h2438; // 0x1a0e
	13'h0d08: q0 = 16'h302d; // 0x1a10
	13'h0d09: q0 = 16'h000e; // 0x1a12
	13'h0d0a: q0 = 16'hc07c; // 0x1a14
	13'h0d0b: q0 = 16'h000f; // 0x1a16
	13'h0d0c: q0 = 16'h6718; // 0x1a18
	13'h0d0d: q0 = 16'h302d; // 0x1a1a
	13'h0d0e: q0 = 16'h000e; // 0x1a1c
	13'h0d0f: q0 = 16'hc07c; // 0x1a1e
	13'h0d10: q0 = 16'h000f; // 0x1a20
	13'h0d11: q0 = 16'hb07c; // 0x1a22
	13'h0d12: q0 = 16'h0001; // 0x1a24
	13'h0d13: q0 = 16'h670a; // 0x1a26
	13'h0d14: q0 = 16'h082d; // 0x1a28
	13'h0d15: q0 = 16'h0005; // 0x1a2a
	13'h0d16: q0 = 16'h000f; // 0x1a2c
	13'h0d17: q0 = 16'h6700; // 0x1a2e
	13'h0d18: q0 = 16'h03be; // 0x1a30
	13'h0d19: q0 = 16'h302d; // 0x1a32
	13'h0d1a: q0 = 16'h000e; // 0x1a34
	13'h0d1b: q0 = 16'hc07c; // 0x1a36
	13'h0d1c: q0 = 16'h000f; // 0x1a38
	13'h0d1d: q0 = 16'h6600; // 0x1a3a
	13'h0d1e: q0 = 16'h009c; // 0x1a3c
	13'h0d1f: q0 = 16'h082d; // 0x1a3e
	13'h0d20: q0 = 16'h0004; // 0x1a40
	13'h0d21: q0 = 16'h000f; // 0x1a42
	13'h0d22: q0 = 16'h6600; // 0x1a44
	13'h0d23: q0 = 16'h0092; // 0x1a46
	13'h0d24: q0 = 16'h082d; // 0x1a48
	13'h0d25: q0 = 16'h0005; // 0x1a4a
	13'h0d26: q0 = 16'h000f; // 0x1a4c
	13'h0d27: q0 = 16'h6600; // 0x1a4e
	13'h0d28: q0 = 16'h0088; // 0x1a50
	13'h0d29: q0 = 16'h4a6d; // 0x1a52
	13'h0d2a: q0 = 16'h0016; // 0x1a54
	13'h0d2b: q0 = 16'h6600; // 0x1a56
	13'h0d2c: q0 = 16'h007c; // 0x1a58
	13'h0d2d: q0 = 16'h206d; // 0x1a5a
	13'h0d2e: q0 = 16'h001e; // 0x1a5c
	13'h0d2f: q0 = 16'h3ea8; // 0x1a5e
	13'h0d30: q0 = 16'h0002; // 0x1a60
	13'h0d31: q0 = 16'h206d; // 0x1a62
	13'h0d32: q0 = 16'h001e; // 0x1a64
	13'h0d33: q0 = 16'h3f10; // 0x1a66
	13'h0d34: q0 = 16'h206d; // 0x1a68
	13'h0d35: q0 = 16'h001a; // 0x1a6a
	13'h0d36: q0 = 16'h3f10; // 0x1a6c
	13'h0d37: q0 = 16'h4eb9; // 0x1a6e
	13'h0d38: q0 = 16'h0000; // 0x1a70
	13'h0d39: q0 = 16'h2b16; // 0x1a72
	13'h0d3a: q0 = 16'h4a9f; // 0x1a74
	13'h0d3b: q0 = 16'h3a80; // 0x1a76
	13'h0d3c: q0 = 16'h3ead; // 0x1a78
	13'h0d3d: q0 = 16'h0002; // 0x1a7a
	13'h0d3e: q0 = 16'h3f15; // 0x1a7c
	13'h0d3f: q0 = 16'h4eb9; // 0x1a7e
	13'h0d40: q0 = 16'h0000; // 0x1a80
	13'h0d41: q0 = 16'h1280; // 0x1a82
	13'h0d42: q0 = 16'h4a5f; // 0x1a84
	13'h0d43: q0 = 16'h3b40; // 0x1a86
	13'h0d44: q0 = 16'h0004; // 0x1a88
	13'h0d45: q0 = 16'h3ead; // 0x1a8a
	13'h0d46: q0 = 16'h0002; // 0x1a8c
	13'h0d47: q0 = 16'h3f15; // 0x1a8e
	13'h0d48: q0 = 16'h4eb9; // 0x1a90
	13'h0d49: q0 = 16'h0000; // 0x1a92
	13'h0d4a: q0 = 16'ha730; // 0x1a94
	13'h0d4b: q0 = 16'h4a5f; // 0x1a96
	13'h0d4c: q0 = 16'h3b40; // 0x1a98
	13'h0d4d: q0 = 16'h0006; // 0x1a9a
	13'h0d4e: q0 = 16'h7020; // 0x1a9c
	13'h0d4f: q0 = 16'h2279; // 0x1a9e
	13'h0d50: q0 = 16'h0001; // 0x1aa0
	13'h0d51: q0 = 16'h7fb8; // 0x1aa2
	13'h0d52: q0 = 16'h3211; // 0x1aa4
	13'h0d53: q0 = 16'he341; // 0x1aa6
	13'h0d54: q0 = 16'h9041; // 0x1aa8
	13'h0d55: q0 = 16'h3d40; // 0x1aaa
	13'h0d56: q0 = 16'hfffc; // 0x1aac
	13'h0d57: q0 = 16'h0c6e; // 0x1aae
	13'h0d58: q0 = 16'h0003; // 0x1ab0
	13'h0d59: q0 = 16'hfffc; // 0x1ab2
	13'h0d5a: q0 = 16'h6e08; // 0x1ab4
	13'h0d5b: q0 = 16'h3b7c; // 0x1ab6
	13'h0d5c: q0 = 16'h0003; // 0x1ab8
	13'h0d5d: q0 = 16'h0016; // 0x1aba
	13'h0d5e: q0 = 16'h6014; // 0x1abc
	13'h0d5f: q0 = 16'h3eae; // 0x1abe
	13'h0d60: q0 = 16'hfffc; // 0x1ac0
	13'h0d61: q0 = 16'h3f3c; // 0x1ac2
	13'h0d62: q0 = 16'h0003; // 0x1ac4
	13'h0d63: q0 = 16'h4eb9; // 0x1ac6
	13'h0d64: q0 = 16'h0000; // 0x1ac8
	13'h0d65: q0 = 16'h8e6c; // 0x1aca
	13'h0d66: q0 = 16'h4a5f; // 0x1acc
	13'h0d67: q0 = 16'h3b40; // 0x1ace
	13'h0d68: q0 = 16'h0016; // 0x1ad0
	13'h0d69: q0 = 16'h6004; // 0x1ad2
	13'h0d6a: q0 = 16'h536d; // 0x1ad4
	13'h0d6b: q0 = 16'h0016; // 0x1ad6
	13'h0d6c: q0 = 16'h082d; // 0x1ad8
	13'h0d6d: q0 = 16'h0000; // 0x1ada
	13'h0d6e: q0 = 16'h000e; // 0x1adc
	13'h0d6f: q0 = 16'h6622; // 0x1ade
	13'h0d70: q0 = 16'h4a6d; // 0x1ae0
	13'h0d71: q0 = 16'h000a; // 0x1ae2
	13'h0d72: q0 = 16'h6618; // 0x1ae4
	13'h0d73: q0 = 16'h3b6d; // 0x1ae6
	13'h0d74: q0 = 16'h000c; // 0x1ae8
	13'h0d75: q0 = 16'h000a; // 0x1aea
	13'h0d76: q0 = 16'h526d; // 0x1aec
	13'h0d77: q0 = 16'h0008; // 0x1aee
	13'h0d78: q0 = 16'h0c6d; // 0x1af0
	13'h0d79: q0 = 16'h0004; // 0x1af2
	13'h0d7a: q0 = 16'h0008; // 0x1af4
	13'h0d7b: q0 = 16'h6d04; // 0x1af6
	13'h0d7c: q0 = 16'h426d; // 0x1af8
	13'h0d7d: q0 = 16'h0008; // 0x1afa
	13'h0d7e: q0 = 16'h6004; // 0x1afc
	13'h0d7f: q0 = 16'h536d; // 0x1afe
	13'h0d80: q0 = 16'h000a; // 0x1b00
	13'h0d81: q0 = 16'h082d; // 0x1b02
	13'h0d82: q0 = 16'h0000; // 0x1b04
	13'h0d83: q0 = 16'h000e; // 0x1b06
	13'h0d84: q0 = 16'h674c; // 0x1b08
	13'h0d85: q0 = 16'h302d; // 0x1b0a
	13'h0d86: q0 = 16'h000c; // 0x1b0c
	13'h0d87: q0 = 16'hd16d; // 0x1b0e
	13'h0d88: q0 = 16'h0008; // 0x1b10
	13'h0d89: q0 = 16'h0c6d; // 0x1b12
	13'h0d8a: q0 = 16'h0047; // 0x1b14
	13'h0d8b: q0 = 16'h0008; // 0x1b16
	13'h0d8c: q0 = 16'h6f06; // 0x1b18
	13'h0d8d: q0 = 16'h046d; // 0x1b1a
	13'h0d8e: q0 = 16'h0048; // 0x1b1c
	13'h0d8f: q0 = 16'h0008; // 0x1b1e
	13'h0d90: q0 = 16'h206d; // 0x1b20
	13'h0d91: q0 = 16'h0022; // 0x1b22
	13'h0d92: q0 = 16'h322d; // 0x1b24
	13'h0d93: q0 = 16'h0008; // 0x1b26
	13'h0d94: q0 = 16'h48c1; // 0x1b28
	13'h0d95: q0 = 16'hd2bc; // 0x1b2a
	13'h0d96: q0 = 16'h0000; // 0x1b2c
	13'h0d97: q0 = 16'hca18; // 0x1b2e
	13'h0d98: q0 = 16'h2241; // 0x1b30
	13'h0d99: q0 = 16'h1211; // 0x1b32
	13'h0d9a: q0 = 16'h4881; // 0x1b34
	13'h0d9b: q0 = 16'hd27c; // 0x1b36
	13'h0d9c: q0 = 16'h005a; // 0x1b38
	13'h0d9d: q0 = 16'h3141; // 0x1b3a
	13'h0d9e: q0 = 16'h0004; // 0x1b3c
	13'h0d9f: q0 = 16'h3ead; // 0x1b3e
	13'h0da0: q0 = 16'h0008; // 0x1b40
	13'h0da1: q0 = 16'h202d; // 0x1b42
	13'h0da2: q0 = 16'h0022; // 0x1b44
	13'h0da3: q0 = 16'h5c80; // 0x1b46
	13'h0da4: q0 = 16'h2f00; // 0x1b48
	13'h0da5: q0 = 16'h4eb9; // 0x1b4a
	13'h0da6: q0 = 16'h0000; // 0x1b4c
	13'h0da7: q0 = 16'h3ee6; // 0x1b4e
	13'h0da8: q0 = 16'h4a9f; // 0x1b50
	13'h0da9: q0 = 16'h6000; // 0x1b52
	13'h0daa: q0 = 16'h00c0; // 0x1b54
	13'h0dab: q0 = 16'h082d; // 0x1b56
	13'h0dac: q0 = 16'h0001; // 0x1b58
	13'h0dad: q0 = 16'h000e; // 0x1b5a
	13'h0dae: q0 = 16'h6600; // 0x1b5c
	13'h0daf: q0 = 16'h00b6; // 0x1b5e
	13'h0db0: q0 = 16'h082d; // 0x1b60
	13'h0db1: q0 = 16'h0004; // 0x1b62
	13'h0db2: q0 = 16'h000f; // 0x1b64
	13'h0db3: q0 = 16'h6712; // 0x1b66
	13'h0db4: q0 = 16'h206d; // 0x1b68
	13'h0db5: q0 = 16'h001e; // 0x1b6a
	13'h0db6: q0 = 16'h322d; // 0x1b6c
	13'h0db7: q0 = 16'h0008; // 0x1b6e
	13'h0db8: q0 = 16'hd27c; // 0x1b70
	13'h0db9: q0 = 16'h00db; // 0x1b72
	13'h0dba: q0 = 16'h3141; // 0x1b74
	13'h0dbb: q0 = 16'h0004; // 0x1b76
	13'h0dbc: q0 = 16'h6028; // 0x1b78
	13'h0dbd: q0 = 16'h4aad; // 0x1b7a
	13'h0dbe: q0 = 16'h0010; // 0x1b7c
	13'h0dbf: q0 = 16'h6612; // 0x1b7e
	13'h0dc0: q0 = 16'h206d; // 0x1b80
	13'h0dc1: q0 = 16'h001e; // 0x1b82
	13'h0dc2: q0 = 16'h322d; // 0x1b84
	13'h0dc3: q0 = 16'h0008; // 0x1b86
	13'h0dc4: q0 = 16'hd27c; // 0x1b88
	13'h0dc5: q0 = 16'h0067; // 0x1b8a
	13'h0dc6: q0 = 16'h3141; // 0x1b8c
	13'h0dc7: q0 = 16'h0004; // 0x1b8e
	13'h0dc8: q0 = 16'h6010; // 0x1b90
	13'h0dc9: q0 = 16'h206d; // 0x1b92
	13'h0dca: q0 = 16'h001e; // 0x1b94
	13'h0dcb: q0 = 16'h322d; // 0x1b96
	13'h0dcc: q0 = 16'h0008; // 0x1b98
	13'h0dcd: q0 = 16'hd27c; // 0x1b9a
	13'h0dce: q0 = 16'h006b; // 0x1b9c
	13'h0dcf: q0 = 16'h3141; // 0x1b9e
	13'h0dd0: q0 = 16'h0004; // 0x1ba0
	13'h0dd1: q0 = 16'h3e95; // 0x1ba2
	13'h0dd2: q0 = 16'h202d; // 0x1ba4
	13'h0dd3: q0 = 16'h001e; // 0x1ba6
	13'h0dd4: q0 = 16'h5c80; // 0x1ba8
	13'h0dd5: q0 = 16'h2f00; // 0x1baa
	13'h0dd6: q0 = 16'h4eb9; // 0x1bac
	13'h0dd7: q0 = 16'h0000; // 0x1bae
	13'h0dd8: q0 = 16'h3ee6; // 0x1bb0
	13'h0dd9: q0 = 16'h4a9f; // 0x1bb2
	13'h0dda: q0 = 16'h082d; // 0x1bb4
	13'h0ddb: q0 = 16'h0004; // 0x1bb6
	13'h0ddc: q0 = 16'h000f; // 0x1bb8
	13'h0ddd: q0 = 16'h671c; // 0x1bba
	13'h0dde: q0 = 16'h206d; // 0x1bbc
	13'h0ddf: q0 = 16'h0022; // 0x1bbe
	13'h0de0: q0 = 16'h322d; // 0x1bc0
	13'h0de1: q0 = 16'h0008; // 0x1bc2
	13'h0de2: q0 = 16'h48c1; // 0x1bc4
	13'h0de3: q0 = 16'hd2bc; // 0x1bc6
	13'h0de4: q0 = 16'h0000; // 0x1bc8
	13'h0de5: q0 = 16'hc880; // 0x1bca
	13'h0de6: q0 = 16'h2241; // 0x1bcc
	13'h0de7: q0 = 16'h1211; // 0x1bce
	13'h0de8: q0 = 16'h4881; // 0x1bd0
	13'h0de9: q0 = 16'h3141; // 0x1bd2
	13'h0dea: q0 = 16'h0004; // 0x1bd4
	13'h0deb: q0 = 16'h602a; // 0x1bd6
	13'h0dec: q0 = 16'h302d; // 0x1bd8
	13'h0ded: q0 = 16'h000e; // 0x1bda
	13'h0dee: q0 = 16'hc07c; // 0x1bdc
	13'h0def: q0 = 16'h000f; // 0x1bde
	13'h0df0: q0 = 16'hb07c; // 0x1be0
	13'h0df1: q0 = 16'h0001; // 0x1be2
	13'h0df2: q0 = 16'h671c; // 0x1be4
	13'h0df3: q0 = 16'h206d; // 0x1be6
	13'h0df4: q0 = 16'h0022; // 0x1be8
	13'h0df5: q0 = 16'h3215; // 0x1bea
	13'h0df6: q0 = 16'h48c1; // 0x1bec
	13'h0df7: q0 = 16'hd2bc; // 0x1bee
	13'h0df8: q0 = 16'h0000; // 0x1bf0
	13'h0df9: q0 = 16'hca18; // 0x1bf2
	13'h0dfa: q0 = 16'h2241; // 0x1bf4
	13'h0dfb: q0 = 16'h1211; // 0x1bf6
	13'h0dfc: q0 = 16'h4881; // 0x1bf8
	13'h0dfd: q0 = 16'hd27c; // 0x1bfa
	13'h0dfe: q0 = 16'h005a; // 0x1bfc
	13'h0dff: q0 = 16'h3141; // 0x1bfe
	13'h0e00: q0 = 16'h0004; // 0x1c00
	13'h0e01: q0 = 16'h3e95; // 0x1c02
	13'h0e02: q0 = 16'h202d; // 0x1c04
	13'h0e03: q0 = 16'h0022; // 0x1c06
	13'h0e04: q0 = 16'h5c80; // 0x1c08
	13'h0e05: q0 = 16'h2f00; // 0x1c0a
	13'h0e06: q0 = 16'h4eb9; // 0x1c0c
	13'h0e07: q0 = 16'h0000; // 0x1c0e
	13'h0e08: q0 = 16'h3ee6; // 0x1c10
	13'h0e09: q0 = 16'h4a9f; // 0x1c12
	13'h0e0a: q0 = 16'h206d; // 0x1c14
	13'h0e0b: q0 = 16'h001e; // 0x1c16
	13'h0e0c: q0 = 16'h3c10; // 0x1c18
	13'h0e0d: q0 = 16'h206d; // 0x1c1a
	13'h0e0e: q0 = 16'h001e; // 0x1c1c
	13'h0e0f: q0 = 16'h3a28; // 0x1c1e
	13'h0e10: q0 = 16'h0002; // 0x1c20
	13'h0e11: q0 = 16'h082d; // 0x1c22
	13'h0e12: q0 = 16'h0004; // 0x1c24
	13'h0e13: q0 = 16'h000f; // 0x1c26
	13'h0e14: q0 = 16'h6718; // 0x1c28
	13'h0e15: q0 = 16'h3a2d; // 0x1c2a
	13'h0e16: q0 = 16'h0008; // 0x1c2c
	13'h0e17: q0 = 16'hef45; // 0x1c2e
	13'h0e18: q0 = 16'hda6d; // 0x1c30
	13'h0e19: q0 = 16'h0018; // 0x1c32
	13'h0e1a: q0 = 16'h0c6d; // 0x1c34
	13'h0e1b: q0 = 16'h0003; // 0x1c36
	13'h0e1c: q0 = 16'h0008; // 0x1c38
	13'h0e1d: q0 = 16'h6604; // 0x1c3a
	13'h0e1e: q0 = 16'h9a7c; // 0x1c3c
	13'h0e1f: q0 = 16'h0100; // 0x1c3e
	13'h0e20: q0 = 16'h6026; // 0x1c40
	13'h0e21: q0 = 16'h082d; // 0x1c42
	13'h0e22: q0 = 16'h0001; // 0x1c44
	13'h0e23: q0 = 16'h000e; // 0x1c46
	13'h0e24: q0 = 16'h671e; // 0x1c48
	13'h0e25: q0 = 16'h3a2d; // 0x1c4a
	13'h0e26: q0 = 16'h0008; // 0x1c4c
	13'h0e27: q0 = 16'hef45; // 0x1c4e
	13'h0e28: q0 = 16'hda6d; // 0x1c50
	13'h0e29: q0 = 16'h0018; // 0x1c52
	13'h0e2a: q0 = 16'h0c6d; // 0x1c54
	13'h0e2b: q0 = 16'h0001; // 0x1c56
	13'h0e2c: q0 = 16'h0008; // 0x1c58
	13'h0e2d: q0 = 16'h6708; // 0x1c5a
	13'h0e2e: q0 = 16'h0c6d; // 0x1c5c
	13'h0e2f: q0 = 16'h0002; // 0x1c5e
	13'h0e30: q0 = 16'h0008; // 0x1c60
	13'h0e31: q0 = 16'h6604; // 0x1c62
	13'h0e32: q0 = 16'hda7c; // 0x1c64
	13'h0e33: q0 = 16'h0100; // 0x1c66
	13'h0e34: q0 = 16'h302d; // 0x1c68
	13'h0e35: q0 = 16'h000e; // 0x1c6a
	13'h0e36: q0 = 16'hc07c; // 0x1c6c
	13'h0e37: q0 = 16'h000f; // 0x1c6e
	13'h0e38: q0 = 16'h6610; // 0x1c70
	13'h0e39: q0 = 16'h082d; // 0x1c72
	13'h0e3a: q0 = 16'h0004; // 0x1c74
	13'h0e3b: q0 = 16'h000f; // 0x1c76
	13'h0e3c: q0 = 16'h6608; // 0x1c78
	13'h0e3d: q0 = 16'h082d; // 0x1c7a
	13'h0e3e: q0 = 16'h0005; // 0x1c7c
	13'h0e3f: q0 = 16'h000f; // 0x1c7e
	13'h0e40: q0 = 16'h6704; // 0x1c80
	13'h0e41: q0 = 16'h4240; // 0x1c82
	13'h0e42: q0 = 16'h6002; // 0x1c84
	13'h0e43: q0 = 16'h7001; // 0x1c86
	13'h0e44: q0 = 16'h3d40; // 0x1c88
	13'h0e45: q0 = 16'hfffe; // 0x1c8a
	13'h0e46: q0 = 16'h302d; // 0x1c8c
	13'h0e47: q0 = 16'h0004; // 0x1c8e
	13'h0e48: q0 = 16'hd046; // 0x1c90
	13'h0e49: q0 = 16'h3c00; // 0x1c92
	13'h0e4a: q0 = 16'hbc7c; // 0x1c94
	13'h0e4b: q0 = 16'h0180; // 0x1c96
	13'h0e4c: q0 = 16'h6c10; // 0x1c98
	13'h0e4d: q0 = 16'h4a6e; // 0x1c9a
	13'h0e4e: q0 = 16'hfffe; // 0x1c9c
	13'h0e4f: q0 = 16'h6706; // 0x1c9e
	13'h0e50: q0 = 16'h3c3c; // 0x1ca0
	13'h0e51: q0 = 16'h0180; // 0x1ca2
	13'h0e52: q0 = 16'h6004; // 0x1ca4
	13'h0e53: q0 = 16'h6000; // 0x1ca6
	13'h0e54: q0 = 16'h013e; // 0x1ca8
	13'h0e55: q0 = 16'hbc7c; // 0x1caa
	13'h0e56: q0 = 16'h7780; // 0x1cac
	13'h0e57: q0 = 16'h6d10; // 0x1cae
	13'h0e58: q0 = 16'h4a6e; // 0x1cb0
	13'h0e59: q0 = 16'hfffe; // 0x1cb2
	13'h0e5a: q0 = 16'h6706; // 0x1cb4
	13'h0e5b: q0 = 16'h3c3c; // 0x1cb6
	13'h0e5c: q0 = 16'h7700; // 0x1cb8
	13'h0e5d: q0 = 16'h6004; // 0x1cba
	13'h0e5e: q0 = 16'h6000; // 0x1cbc
	13'h0e5f: q0 = 16'h0128; // 0x1cbe
	13'h0e60: q0 = 16'h302d; // 0x1cc0
	13'h0e61: q0 = 16'h0006; // 0x1cc2
	13'h0e62: q0 = 16'hd045; // 0x1cc4
	13'h0e63: q0 = 16'h3a00; // 0x1cc6
	13'h0e64: q0 = 16'hba7c; // 0x1cc8
	13'h0e65: q0 = 16'h1400; // 0x1cca
	13'h0e66: q0 = 16'h6c10; // 0x1ccc
	13'h0e67: q0 = 16'h4a6e; // 0x1cce
	13'h0e68: q0 = 16'hfffe; // 0x1cd0
	13'h0e69: q0 = 16'h6706; // 0x1cd2
	13'h0e6a: q0 = 16'h3a3c; // 0x1cd4
	13'h0e6b: q0 = 16'h1400; // 0x1cd6
	13'h0e6c: q0 = 16'h6004; // 0x1cd8
	13'h0e6d: q0 = 16'h6000; // 0x1cda
	13'h0e6e: q0 = 16'h010a; // 0x1cdc
	13'h0e6f: q0 = 16'hba7c; // 0x1cde
	13'h0e70: q0 = 16'h7400; // 0x1ce0
	13'h0e71: q0 = 16'h6d18; // 0x1ce2
	13'h0e72: q0 = 16'h082d; // 0x1ce4
	13'h0e73: q0 = 16'h0004; // 0x1ce6
	13'h0e74: q0 = 16'h000f; // 0x1ce8
	13'h0e75: q0 = 16'h6610; // 0x1cea
	13'h0e76: q0 = 16'h4a6e; // 0x1cec
	13'h0e77: q0 = 16'hfffe; // 0x1cee
	13'h0e78: q0 = 16'h6706; // 0x1cf0
	13'h0e79: q0 = 16'h3a3c; // 0x1cf2
	13'h0e7a: q0 = 16'h7380; // 0x1cf4
	13'h0e7b: q0 = 16'h6004; // 0x1cf6
	13'h0e7c: q0 = 16'h6000; // 0x1cf8
	13'h0e7d: q0 = 16'h00ec; // 0x1cfa
	13'h0e7e: q0 = 16'h082d; // 0x1cfc
	13'h0e7f: q0 = 16'h0004; // 0x1cfe
	13'h0e80: q0 = 16'h000f; // 0x1d00
	13'h0e81: q0 = 16'h6604; // 0x1d02
	13'h0e82: q0 = 16'h3b45; // 0x1d04
	13'h0e83: q0 = 16'h0018; // 0x1d06
	13'h0e84: q0 = 16'h3e85; // 0x1d08
	13'h0e85: q0 = 16'h3f06; // 0x1d0a
	13'h0e86: q0 = 16'h2f0d; // 0x1d0c
	13'h0e87: q0 = 16'h4eb9; // 0x1d0e
	13'h0e88: q0 = 16'h0000; // 0x1d10
	13'h0e89: q0 = 16'h2dc2; // 0x1d12
	13'h0e8a: q0 = 16'h5c4f; // 0x1d14
	13'h0e8b: q0 = 16'h4aad; // 0x1d16
	13'h0e8c: q0 = 16'h0010; // 0x1d18
	13'h0e8d: q0 = 16'h6742; // 0x1d1a
	13'h0e8e: q0 = 16'h0c55; // 0x1d1c
	13'h0e8f: q0 = 16'h0012; // 0x1d1e
	13'h0e90: q0 = 16'h6f12; // 0x1d20
	13'h0e91: q0 = 16'h0c55; // 0x1d22
	13'h0e92: q0 = 16'h0036; // 0x1d24
	13'h0e93: q0 = 16'h6e0c; // 0x1d26
	13'h0e94: q0 = 16'h206d; // 0x1d28
	13'h0e95: q0 = 16'h001e; // 0x1d2a
	13'h0e96: q0 = 16'h3c10; // 0x1d2c
	13'h0e97: q0 = 16'hdc7c; // 0x1d2e
	13'h0e98: q0 = 16'h0280; // 0x1d30
	13'h0e99: q0 = 16'h600a; // 0x1d32
	13'h0e9a: q0 = 16'h206d; // 0x1d34
	13'h0e9b: q0 = 16'h001e; // 0x1d36
	13'h0e9c: q0 = 16'h3c10; // 0x1d38
	13'h0e9d: q0 = 16'hdc7c; // 0x1d3a
	13'h0e9e: q0 = 16'hfd80; // 0x1d3c
	13'h0e9f: q0 = 16'h206d; // 0x1d3e
	13'h0ea0: q0 = 16'h001e; // 0x1d40
	13'h0ea1: q0 = 16'h3a28; // 0x1d42
	13'h0ea2: q0 = 16'h0002; // 0x1d44
	13'h0ea3: q0 = 16'hda7c; // 0x1d46
	13'h0ea4: q0 = 16'h0180; // 0x1d48
	13'h0ea5: q0 = 16'h3ebc; // 0x1d4a
	13'h0ea6: q0 = 16'h0001; // 0x1d4c
	13'h0ea7: q0 = 16'h3f05; // 0x1d4e
	13'h0ea8: q0 = 16'h3f06; // 0x1d50
	13'h0ea9: q0 = 16'h2f2d; // 0x1d52
	13'h0eaa: q0 = 16'h0010; // 0x1d54
	13'h0eab: q0 = 16'h4eb9; // 0x1d56
	13'h0eac: q0 = 16'h0000; // 0x1d58
	13'h0ead: q0 = 16'h3c92; // 0x1d5a
	13'h0eae: q0 = 16'hbf8f; // 0x1d5c
	13'h0eaf: q0 = 16'h2079; // 0x1d5e
	13'h0eb0: q0 = 16'h0001; // 0x1d60
	13'h0eb1: q0 = 16'h7fb8; // 0x1d62
	13'h0eb2: q0 = 16'h0c50; // 0x1d64
	13'h0eb3: q0 = 16'h0002; // 0x1d66
	13'h0eb4: q0 = 16'h6d00; // 0x1d68
	13'h0eb5: q0 = 16'h0084; // 0x1d6a
	13'h0eb6: q0 = 16'h082d; // 0x1d6c
	13'h0eb7: q0 = 16'h0005; // 0x1d6e
	13'h0eb8: q0 = 16'h000f; // 0x1d70
	13'h0eb9: q0 = 16'h6600; // 0x1d72
	13'h0eba: q0 = 16'h007a; // 0x1d74
	13'h0ebb: q0 = 16'h082d; // 0x1d76
	13'h0ebc: q0 = 16'h0004; // 0x1d78
	13'h0ebd: q0 = 16'h000f; // 0x1d7a
	13'h0ebe: q0 = 16'h6600; // 0x1d7c
	13'h0ebf: q0 = 16'h0070; // 0x1d7e
	13'h0ec0: q0 = 16'h302d; // 0x1d80
	13'h0ec1: q0 = 16'h000e; // 0x1d82
	13'h0ec2: q0 = 16'hc07c; // 0x1d84
	13'h0ec3: q0 = 16'h000f; // 0x1d86
	13'h0ec4: q0 = 16'h6664; // 0x1d88
	13'h0ec5: q0 = 16'h4aad; // 0x1d8a
	13'h0ec6: q0 = 16'h0010; // 0x1d8c
	13'h0ec7: q0 = 16'h663a; // 0x1d8e
	13'h0ec8: q0 = 16'h3ebc; // 0x1d90
	13'h0ec9: q0 = 16'h0001; // 0x1d92
	13'h0eca: q0 = 16'h206d; // 0x1d94
	13'h0ecb: q0 = 16'h001e; // 0x1d96
	13'h0ecc: q0 = 16'h3f28; // 0x1d98
	13'h0ecd: q0 = 16'h0002; // 0x1d9a
	13'h0ece: q0 = 16'h206d; // 0x1d9c
	13'h0ecf: q0 = 16'h001e; // 0x1d9e
	13'h0ed0: q0 = 16'h3f10; // 0x1da0
	13'h0ed1: q0 = 16'h4eb9; // 0x1da2
	13'h0ed2: q0 = 16'h0000; // 0x1da4
	13'h0ed3: q0 = 16'h37e6; // 0x1da6
	13'h0ed4: q0 = 16'h4a9f; // 0x1da8
	13'h0ed5: q0 = 16'h2b40; // 0x1daa
	13'h0ed6: q0 = 16'h0010; // 0x1dac
	13'h0ed7: q0 = 16'h4aad; // 0x1dae
	13'h0ed8: q0 = 16'h0010; // 0x1db0
	13'h0ed9: q0 = 16'h670a; // 0x1db2
	13'h0eda: q0 = 16'h3079; // 0x1db4
	13'h0edb: q0 = 16'h0001; // 0x1db6
	13'h0edc: q0 = 16'h7f28; // 0x1db8
	13'h0edd: q0 = 16'h2b48; // 0x1dba
	13'h0ede: q0 = 16'h002a; // 0x1dbc
	13'h0edf: q0 = 16'h4aad; // 0x1dbe
	13'h0ee0: q0 = 16'h002a; // 0x1dc0
	13'h0ee1: q0 = 16'h6c04; // 0x1dc2
	13'h0ee2: q0 = 16'h42ad; // 0x1dc4
	13'h0ee3: q0 = 16'h002a; // 0x1dc6
	13'h0ee4: q0 = 16'h601a; // 0x1dc8
	13'h0ee5: q0 = 16'h4aad; // 0x1dca
	13'h0ee6: q0 = 16'h002a; // 0x1dcc
	13'h0ee7: q0 = 16'h6614; // 0x1dce
	13'h0ee8: q0 = 16'h2e8d; // 0x1dd0
	13'h0ee9: q0 = 16'h3f15; // 0x1dd2
	13'h0eea: q0 = 16'h2f2d; // 0x1dd4
	13'h0eeb: q0 = 16'h0010; // 0x1dd6
	13'h0eec: q0 = 16'h4eb9; // 0x1dd8
	13'h0eed: q0 = 16'h0000; // 0x1dda
	13'h0eee: q0 = 16'h3b8e; // 0x1ddc
	13'h0eef: q0 = 16'h5c4f; // 0x1dde
	13'h0ef0: q0 = 16'h42ad; // 0x1de0
	13'h0ef1: q0 = 16'h0010; // 0x1de2
	13'h0ef2: q0 = 16'h6008; // 0x1de4
	13'h0ef3: q0 = 16'h2e8d; // 0x1de6
	13'h0ef4: q0 = 16'h4eb9; // 0x1de8
	13'h0ef5: q0 = 16'h0000; // 0x1dea
	13'h0ef6: q0 = 16'h2ec2; // 0x1dec
	13'h0ef7: q0 = 16'hdbfc; // 0x1dee
	13'h0ef8: q0 = 16'h0000; // 0x1df0
	13'h0ef9: q0 = 16'h002e; // 0x1df2
	13'h0efa: q0 = 16'h5247; // 0x1df4
	13'h0efb: q0 = 16'h6000; // 0x1df6
	13'h0efc: q0 = 16'hfb0c; // 0x1df8
	13'h0efd: q0 = 16'h4a9f; // 0x1dfa
	13'h0efe: q0 = 16'h4cdf; // 0x1dfc
	13'h0eff: q0 = 16'h20e0; // 0x1dfe
	13'h0f00: q0 = 16'h4e5e; // 0x1e00
	13'h0f01: q0 = 16'h4e75; // 0x1e02
	13'h0f02: q0 = 16'h4e56; // 0x1e04
	13'h0f03: q0 = 16'h0000; // 0x1e06
	13'h0f04: q0 = 16'h48e7; // 0x1e08
	13'h0f05: q0 = 16'h0f04; // 0x1e0a
	13'h0f06: q0 = 16'h2a7c; // 0x1e0c
	13'h0f07: q0 = 16'h0001; // 0x1e0e
	13'h0f08: q0 = 16'h89be; // 0x1e10
	13'h0f09: q0 = 16'h4247; // 0x1e12
	13'h0f0a: q0 = 16'hbe79; // 0x1e14
	13'h0f0b: q0 = 16'h0001; // 0x1e16
	13'h0f0c: q0 = 16'h7fbc; // 0x1e18
	13'h0f0d: q0 = 16'h6c62; // 0x1e1a
	13'h0f0e: q0 = 16'h302d; // 0x1e1c
	13'h0f0f: q0 = 16'h000e; // 0x1e1e
	13'h0f10: q0 = 16'hc07c; // 0x1e20
	13'h0f11: q0 = 16'h000f; // 0x1e22
	13'h0f12: q0 = 16'h664e; // 0x1e24
	13'h0f13: q0 = 16'h3eae; // 0x1e26
	13'h0f14: q0 = 16'h0008; // 0x1e28
	13'h0f15: q0 = 16'h206d; // 0x1e2a
	13'h0f16: q0 = 16'h001e; // 0x1e2c
	13'h0f17: q0 = 16'h3010; // 0x1e2e
	13'h0f18: q0 = 16'h9157; // 0x1e30
	13'h0f19: q0 = 16'h4eb9; // 0x1e32
	13'h0f1a: q0 = 16'h0000; // 0x1e34
	13'h0f1b: q0 = 16'h09a2; // 0x1e36
	13'h0f1c: q0 = 16'h3c00; // 0x1e38
	13'h0f1d: q0 = 16'h3eae; // 0x1e3a
	13'h0f1e: q0 = 16'h000a; // 0x1e3c
	13'h0f1f: q0 = 16'h206d; // 0x1e3e
	13'h0f20: q0 = 16'h001e; // 0x1e40
	13'h0f21: q0 = 16'h3028; // 0x1e42
	13'h0f22: q0 = 16'h0002; // 0x1e44
	13'h0f23: q0 = 16'h9157; // 0x1e46
	13'h0f24: q0 = 16'h4eb9; // 0x1e48
	13'h0f25: q0 = 16'h0000; // 0x1e4a
	13'h0f26: q0 = 16'h09a2; // 0x1e4c
	13'h0f27: q0 = 16'h3a00; // 0x1e4e
	13'h0f28: q0 = 16'hbc7c; // 0x1e50
	13'h0f29: q0 = 16'h0a00; // 0x1e52
	13'h0f2a: q0 = 16'h6c0c; // 0x1e54
	13'h0f2b: q0 = 16'hba7c; // 0x1e56
	13'h0f2c: q0 = 16'h0a00; // 0x1e58
	13'h0f2d: q0 = 16'h6c06; // 0x1e5a
	13'h0f2e: q0 = 16'h5279; // 0x1e5c
	13'h0f2f: q0 = 16'h0001; // 0x1e5e
	13'h0f30: q0 = 16'h7efc; // 0x1e60
	13'h0f31: q0 = 16'hbc7c; // 0x1e62
	13'h0f32: q0 = 16'h0400; // 0x1e64
	13'h0f33: q0 = 16'h6c0c; // 0x1e66
	13'h0f34: q0 = 16'hba7c; // 0x1e68
	13'h0f35: q0 = 16'h0400; // 0x1e6a
	13'h0f36: q0 = 16'h6c06; // 0x1e6c
	13'h0f37: q0 = 16'h3007; // 0x1e6e
	13'h0f38: q0 = 16'h5240; // 0x1e70
	13'h0f39: q0 = 16'h600c; // 0x1e72
	13'h0f3a: q0 = 16'hdbfc; // 0x1e74
	13'h0f3b: q0 = 16'h0000; // 0x1e76
	13'h0f3c: q0 = 16'h002e; // 0x1e78
	13'h0f3d: q0 = 16'h5247; // 0x1e7a
	13'h0f3e: q0 = 16'h6096; // 0x1e7c
	13'h0f3f: q0 = 16'h4240; // 0x1e7e
	13'h0f40: q0 = 16'h4a9f; // 0x1e80
	13'h0f41: q0 = 16'h4cdf; // 0x1e82
	13'h0f42: q0 = 16'h20e0; // 0x1e84
	13'h0f43: q0 = 16'h4e5e; // 0x1e86
	13'h0f44: q0 = 16'h4e75; // 0x1e88
	13'h0f45: q0 = 16'h4e56; // 0x1e8a
	13'h0f46: q0 = 16'h0000; // 0x1e8c
	13'h0f47: q0 = 16'h48e7; // 0x1e8e
	13'h0f48: q0 = 16'h0304; // 0x1e90
	13'h0f49: q0 = 16'h2a7c; // 0x1e92
	13'h0f4a: q0 = 16'h0001; // 0x1e94
	13'h0f4b: q0 = 16'h89be; // 0x1e96
	13'h0f4c: q0 = 16'h4247; // 0x1e98
	13'h0f4d: q0 = 16'hbe7c; // 0x1e9a
	13'h0f4e: q0 = 16'h0004; // 0x1e9c
	13'h0f4f: q0 = 16'h6c6a; // 0x1e9e
	13'h0f50: q0 = 16'h206d; // 0x1ea0
	13'h0f51: q0 = 16'h001e; // 0x1ea2
	13'h0f52: q0 = 16'h317c; // 0x1ea4
	13'h0f53: q0 = 16'h0030; // 0x1ea6
	13'h0f54: q0 = 16'h0004; // 0x1ea8
	13'h0f55: q0 = 16'h206d; // 0x1eaa
	13'h0f56: q0 = 16'h0022; // 0x1eac
	13'h0f57: q0 = 16'h317c; // 0x1eae
	13'h0f58: q0 = 16'h0030; // 0x1eb0
	13'h0f59: q0 = 16'h0004; // 0x1eb2
	13'h0f5a: q0 = 16'h206d; // 0x1eb4
	13'h0f5b: q0 = 16'h0026; // 0x1eb6
	13'h0f5c: q0 = 16'h317c; // 0x1eb8
	13'h0f5d: q0 = 16'h0030; // 0x1eba
	13'h0f5e: q0 = 16'h0004; // 0x1ebc
	13'h0f5f: q0 = 16'h206d; // 0x1ebe
	13'h0f60: q0 = 16'h001e; // 0x1ec0
	13'h0f61: q0 = 16'h4250; // 0x1ec2
	13'h0f62: q0 = 16'h206d; // 0x1ec4
	13'h0f63: q0 = 16'h001e; // 0x1ec6
	13'h0f64: q0 = 16'h4268; // 0x1ec8
	13'h0f65: q0 = 16'h0002; // 0x1eca
	13'h0f66: q0 = 16'h206d; // 0x1ecc
	13'h0f67: q0 = 16'h001e; // 0x1ece
	13'h0f68: q0 = 16'h4268; // 0x1ed0
	13'h0f69: q0 = 16'h0006; // 0x1ed2
	13'h0f6a: q0 = 16'h206d; // 0x1ed4
	13'h0f6b: q0 = 16'h0022; // 0x1ed6
	13'h0f6c: q0 = 16'h4250; // 0x1ed8
	13'h0f6d: q0 = 16'h206d; // 0x1eda
	13'h0f6e: q0 = 16'h0022; // 0x1edc
	13'h0f6f: q0 = 16'h4268; // 0x1ede
	13'h0f70: q0 = 16'h0002; // 0x1ee0
	13'h0f71: q0 = 16'h206d; // 0x1ee2
	13'h0f72: q0 = 16'h0022; // 0x1ee4
	13'h0f73: q0 = 16'h4268; // 0x1ee6
	13'h0f74: q0 = 16'h0006; // 0x1ee8
	13'h0f75: q0 = 16'h206d; // 0x1eea
	13'h0f76: q0 = 16'h0026; // 0x1eec
	13'h0f77: q0 = 16'h4250; // 0x1eee
	13'h0f78: q0 = 16'h206d; // 0x1ef0
	13'h0f79: q0 = 16'h0026; // 0x1ef2
	13'h0f7a: q0 = 16'h4268; // 0x1ef4
	13'h0f7b: q0 = 16'h0002; // 0x1ef6
	13'h0f7c: q0 = 16'h206d; // 0x1ef8
	13'h0f7d: q0 = 16'h0026; // 0x1efa
	13'h0f7e: q0 = 16'h4268; // 0x1efc
	13'h0f7f: q0 = 16'h0006; // 0x1efe
	13'h0f80: q0 = 16'hdbfc; // 0x1f00
	13'h0f81: q0 = 16'h0000; // 0x1f02
	13'h0f82: q0 = 16'h002e; // 0x1f04
	13'h0f83: q0 = 16'h5247; // 0x1f06
	13'h0f84: q0 = 16'h6090; // 0x1f08
	13'h0f85: q0 = 16'h4279; // 0x1f0a
	13'h0f86: q0 = 16'h0001; // 0x1f0c
	13'h0f87: q0 = 16'h86d4; // 0x1f0e
	13'h0f88: q0 = 16'h4a9f; // 0x1f10
	13'h0f89: q0 = 16'h4cdf; // 0x1f12
	13'h0f8a: q0 = 16'h2080; // 0x1f14
	13'h0f8b: q0 = 16'h4e5e; // 0x1f16
	13'h0f8c: q0 = 16'h4e75; // 0x1f18
	13'h0f8d: q0 = 16'h4e56; // 0x1f1a
	13'h0f8e: q0 = 16'h0000; // 0x1f1c
	13'h0f8f: q0 = 16'h48e7; // 0x1f1e
	13'h0f90: q0 = 16'h0104; // 0x1f20
	13'h0f91: q0 = 16'h302e; // 0x1f22
	13'h0f92: q0 = 16'h0008; // 0x1f24
	13'h0f93: q0 = 16'h5340; // 0x1f26
	13'h0f94: q0 = 16'hc1fc; // 0x1f28
	13'h0f95: q0 = 16'h002e; // 0x1f2a
	13'h0f96: q0 = 16'h2a40; // 0x1f2c
	13'h0f97: q0 = 16'hdbfc; // 0x1f2e
	13'h0f98: q0 = 16'h0001; // 0x1f30
	13'h0f99: q0 = 16'h89be; // 0x1f32
	13'h0f9a: q0 = 16'h42ad; // 0x1f34
	13'h0f9b: q0 = 16'h002a; // 0x1f36
	13'h0f9c: q0 = 16'h3eae; // 0x1f38
	13'h0f9d: q0 = 16'h0008; // 0x1f3a
	13'h0f9e: q0 = 16'h2f0d; // 0x1f3c
	13'h0f9f: q0 = 16'h4eb9; // 0x1f3e
	13'h0fa0: q0 = 16'h0000; // 0x1f40
	13'h0fa1: q0 = 16'h2c02; // 0x1f42
	13'h0fa2: q0 = 16'h4a9f; // 0x1f44
	13'h0fa3: q0 = 16'h4a9f; // 0x1f46
	13'h0fa4: q0 = 16'h4cdf; // 0x1f48
	13'h0fa5: q0 = 16'h2000; // 0x1f4a
	13'h0fa6: q0 = 16'h4e5e; // 0x1f4c
	13'h0fa7: q0 = 16'h4e75; // 0x1f4e
	13'h0fa8: q0 = 16'h4e56; // 0x1f50
	13'h0fa9: q0 = 16'h0000; // 0x1f52
	13'h0faa: q0 = 16'h48e7; // 0x1f54
	13'h0fab: q0 = 16'h0104; // 0x1f56
	13'h0fac: q0 = 16'h2a6e; // 0x1f58
	13'h0fad: q0 = 16'h0008; // 0x1f5a
	13'h0fae: q0 = 16'h206d; // 0x1f5c
	13'h0faf: q0 = 16'h001e; // 0x1f5e
	13'h0fb0: q0 = 16'h3ea8; // 0x1f60
	13'h0fb1: q0 = 16'h0002; // 0x1f62
	13'h0fb2: q0 = 16'h206d; // 0x1f64
	13'h0fb3: q0 = 16'h001e; // 0x1f66
	13'h0fb4: q0 = 16'h3f10; // 0x1f68
	13'h0fb5: q0 = 16'h4eb9; // 0x1f6a
	13'h0fb6: q0 = 16'h0000; // 0x1f6c
	13'h0fb7: q0 = 16'h5eb0; // 0x1f6e
	13'h0fb8: q0 = 16'h4a5f; // 0x1f70
	13'h0fb9: q0 = 16'h4eb9; // 0x1f72
	13'h0fba: q0 = 16'h0000; // 0x1f74
	13'h0fbb: q0 = 16'h4738; // 0x1f76
	13'h0fbc: q0 = 16'hb07c; // 0x1f78
	13'h0fbd: q0 = 16'h0002; // 0x1f7a
	13'h0fbe: q0 = 16'h671e; // 0x1f7c
	13'h0fbf: q0 = 16'h206d; // 0x1f7e
	13'h0fc0: q0 = 16'h001e; // 0x1f80
	13'h0fc1: q0 = 16'h317c; // 0x1f82
	13'h0fc2: q0 = 16'h0009; // 0x1f84
	13'h0fc3: q0 = 16'h0006; // 0x1f86
	13'h0fc4: q0 = 16'h206d; // 0x1f88
	13'h0fc5: q0 = 16'h0022; // 0x1f8a
	13'h0fc6: q0 = 16'h317c; // 0x1f8c
	13'h0fc7: q0 = 16'h0008; // 0x1f8e
	13'h0fc8: q0 = 16'h0006; // 0x1f90
	13'h0fc9: q0 = 16'h206d; // 0x1f92
	13'h0fca: q0 = 16'h0026; // 0x1f94
	13'h0fcb: q0 = 16'h317c; // 0x1f96
	13'h0fcc: q0 = 16'h0009; // 0x1f98
	13'h0fcd: q0 = 16'h0006; // 0x1f9a
	13'h0fce: q0 = 16'h206d; // 0x1f9c
	13'h0fcf: q0 = 16'h001e; // 0x1f9e
	13'h0fd0: q0 = 16'h317c; // 0x1fa0
	13'h0fd1: q0 = 16'h0067; // 0x1fa2
	13'h0fd2: q0 = 16'h0004; // 0x1fa4
	13'h0fd3: q0 = 16'h3e95; // 0x1fa6
	13'h0fd4: q0 = 16'h202d; // 0x1fa8
	13'h0fd5: q0 = 16'h001e; // 0x1faa
	13'h0fd6: q0 = 16'h5c80; // 0x1fac
	13'h0fd7: q0 = 16'h2f00; // 0x1fae
	13'h0fd8: q0 = 16'h4eb9; // 0x1fb0
	13'h0fd9: q0 = 16'h0000; // 0x1fb2
	13'h0fda: q0 = 16'h3ee6; // 0x1fb4
	13'h0fdb: q0 = 16'h4a9f; // 0x1fb6
	13'h0fdc: q0 = 16'h3e95; // 0x1fb8
	13'h0fdd: q0 = 16'h202d; // 0x1fba
	13'h0fde: q0 = 16'h0022; // 0x1fbc
	13'h0fdf: q0 = 16'h5c80; // 0x1fbe
	13'h0fe0: q0 = 16'h2f00; // 0x1fc0
	13'h0fe1: q0 = 16'h4eb9; // 0x1fc2
	13'h0fe2: q0 = 16'h0000; // 0x1fc4
	13'h0fe3: q0 = 16'h3ee6; // 0x1fc6
	13'h0fe4: q0 = 16'h4a9f; // 0x1fc8
	13'h0fe5: q0 = 16'h206d; // 0x1fca
	13'h0fe6: q0 = 16'h001a; // 0x1fcc
	13'h0fe7: q0 = 16'h3028; // 0x1fce
	13'h0fe8: q0 = 16'h0002; // 0x1fd0
	13'h0fe9: q0 = 16'h2279; // 0x1fd2
	13'h0fea: q0 = 16'h0001; // 0x1fd4
	13'h0feb: q0 = 16'h7fb8; // 0x1fd6
	13'h0fec: q0 = 16'h3211; // 0x1fd8
	13'h0fed: q0 = 16'h5341; // 0x1fda
	13'h0fee: q0 = 16'he541; // 0x1fdc
	13'h0fef: q0 = 16'hd041; // 0x1fde
	13'h0ff0: q0 = 16'h3b40; // 0x1fe0
	13'h0ff1: q0 = 16'h0002; // 0x1fe2
	13'h0ff2: q0 = 16'h206d; // 0x1fe4
	13'h0ff3: q0 = 16'h001a; // 0x1fe6
	13'h0ff4: q0 = 16'h3028; // 0x1fe8
	13'h0ff5: q0 = 16'h0004; // 0x1fea
	13'h0ff6: q0 = 16'h2279; // 0x1fec
	13'h0ff7: q0 = 16'h0001; // 0x1fee
	13'h0ff8: q0 = 16'h7fb8; // 0x1ff0
	13'h0ff9: q0 = 16'h3211; // 0x1ff2
	13'h0ffa: q0 = 16'he441; // 0x1ff4
	13'h0ffb: q0 = 16'h9041; // 0x1ff6
	13'h0ffc: q0 = 16'h3b40; // 0x1ff8
	13'h0ffd: q0 = 16'h000c; // 0x1ffa
	13'h0ffe: q0 = 16'h4a6d; // 0x1ffc
	13'h0fff: q0 = 16'h000c; // 0x1ffe
	13'h1000: q0 = 16'h6c04; // 0x2000
	13'h1001: q0 = 16'h426d; // 0x2002
	13'h1002: q0 = 16'h000c; // 0x2004
	13'h1003: q0 = 16'h3b6d; // 0x2006
	13'h1004: q0 = 16'h000c; // 0x2008
	13'h1005: q0 = 16'h000a; // 0x200a
	13'h1006: q0 = 16'h426d; // 0x200c
	13'h1007: q0 = 16'h0008; // 0x200e
	13'h1008: q0 = 16'h3b7c; // 0x2010
	13'h1009: q0 = 16'h0010; // 0x2012
	13'h100a: q0 = 16'h0014; // 0x2014
	13'h100b: q0 = 16'h426d; // 0x2016
	13'h100c: q0 = 16'h0016; // 0x2018
	13'h100d: q0 = 16'h426d; // 0x201a
	13'h100e: q0 = 16'h000e; // 0x201c
	13'h100f: q0 = 16'h4a9f; // 0x201e
	13'h1010: q0 = 16'h4cdf; // 0x2020
	13'h1011: q0 = 16'h2000; // 0x2022
	13'h1012: q0 = 16'h4e5e; // 0x2024
	13'h1013: q0 = 16'h4e75; // 0x2026
	13'h1014: q0 = 16'h4e56; // 0x2028
	13'h1015: q0 = 16'h0000; // 0x202a
	13'h1016: q0 = 16'h48e7; // 0x202c
	13'h1017: q0 = 16'h1f04; // 0x202e
	13'h1018: q0 = 16'h2a7c; // 0x2030
	13'h1019: q0 = 16'h0001; // 0x2032
	13'h101a: q0 = 16'h7fde; // 0x2034
	13'h101b: q0 = 16'h4247; // 0x2036
	13'h101c: q0 = 16'h4245; // 0x2038
	13'h101d: q0 = 16'hba7c; // 0x203a
	13'h101e: q0 = 16'h0005; // 0x203c
	13'h101f: q0 = 16'h6c50; // 0x203e
	13'h1020: q0 = 16'h7c01; // 0x2040
	13'h1021: q0 = 16'h4244; // 0x2042
	13'h1022: q0 = 16'h3005; // 0x2044
	13'h1023: q0 = 16'he340; // 0x2046
	13'h1024: q0 = 16'h48c0; // 0x2048
	13'h1025: q0 = 16'hd0bc; // 0x204a
	13'h1026: q0 = 16'h0000; // 0x204c
	13'h1027: q0 = 16'hc7c6; // 0x204e
	13'h1028: q0 = 16'h2040; // 0x2050
	13'h1029: q0 = 16'h3010; // 0x2052
	13'h102a: q0 = 16'hb044; // 0x2054
	13'h102b: q0 = 16'h6f06; // 0x2056
	13'h102c: q0 = 16'hdc5d; // 0x2058
	13'h102d: q0 = 16'h5244; // 0x205a
	13'h102e: q0 = 16'h60e6; // 0x205c
	13'h102f: q0 = 16'h3005; // 0x205e
	13'h1030: q0 = 16'he340; // 0x2060
	13'h1031: q0 = 16'h48c0; // 0x2062
	13'h1032: q0 = 16'hd0bc; // 0x2064
	13'h1033: q0 = 16'h0001; // 0x2066
	13'h1034: q0 = 16'h7fd4; // 0x2068
	13'h1035: q0 = 16'h2040; // 0x206a
	13'h1036: q0 = 16'h3010; // 0x206c
	13'h1037: q0 = 16'hb046; // 0x206e
	13'h1038: q0 = 16'h670a; // 0x2070
	13'h1039: q0 = 16'h7001; // 0x2072
	13'h103a: q0 = 16'h4281; // 0x2074
	13'h103b: q0 = 16'h3205; // 0x2076
	13'h103c: q0 = 16'he360; // 0x2078
	13'h103d: q0 = 16'h8e40; // 0x207a
	13'h103e: q0 = 16'h3005; // 0x207c
	13'h103f: q0 = 16'he340; // 0x207e
	13'h1040: q0 = 16'h48c0; // 0x2080
	13'h1041: q0 = 16'hd0bc; // 0x2082
	13'h1042: q0 = 16'h0001; // 0x2084
	13'h1043: q0 = 16'h7fd4; // 0x2086
	13'h1044: q0 = 16'h2040; // 0x2088
	13'h1045: q0 = 16'h3086; // 0x208a
	13'h1046: q0 = 16'h5245; // 0x208c
	13'h1047: q0 = 16'h60aa; // 0x208e
	13'h1048: q0 = 16'h3007; // 0x2090
	13'h1049: q0 = 16'h4a9f; // 0x2092
	13'h104a: q0 = 16'h4cdf; // 0x2094
	13'h104b: q0 = 16'h20f0; // 0x2096
	13'h104c: q0 = 16'h4e5e; // 0x2098
	13'h104d: q0 = 16'h4e75; // 0x209a
	13'h104e: q0 = 16'h4e56; // 0x209c
	13'h104f: q0 = 16'hffec; // 0x209e
	13'h1050: q0 = 16'h48e7; // 0x20a0
	13'h1051: q0 = 16'h3f1c; // 0x20a2
	13'h1052: q0 = 16'h267c; // 0x20a4
	13'h1053: q0 = 16'h0001; // 0x20a6
	13'h1054: q0 = 16'h7fd4; // 0x20a8
	13'h1055: q0 = 16'h2a79; // 0x20aa
	13'h1056: q0 = 16'h0000; // 0x20ac
	13'h1057: q0 = 16'hc7d0; // 0x20ae
	13'h1058: q0 = 16'h4255; // 0x20b0
	13'h1059: q0 = 16'h287c; // 0x20b2
	13'h105a: q0 = 16'h0001; // 0x20b4
	13'h105b: q0 = 16'h7fd4; // 0x20b6
	13'h105c: q0 = 16'h2a79; // 0x20b8
	13'h105d: q0 = 16'h0000; // 0x20ba
	13'h105e: q0 = 16'hc7d4; // 0x20bc
	13'h105f: q0 = 16'h4246; // 0x20be
	13'h1060: q0 = 16'hbc7c; // 0x20c0
	13'h1061: q0 = 16'h0020; // 0x20c2
	13'h1062: q0 = 16'h6c34; // 0x20c4
	13'h1063: q0 = 16'h301d; // 0x20c6
	13'h1064: q0 = 16'hc07c; // 0x20c8
	13'h1065: q0 = 16'h000f; // 0x20ca
	13'h1066: q0 = 16'h48c0; // 0x20cc
	13'h1067: q0 = 16'h2880; // 0x20ce
	13'h1068: q0 = 16'h7a01; // 0x20d0
	13'h1069: q0 = 16'hba7c; // 0x20d2
	13'h106a: q0 = 16'h0008; // 0x20d4
	13'h106b: q0 = 16'h6c1c; // 0x20d6
	13'h106c: q0 = 16'h3015; // 0x20d8
	13'h106d: q0 = 16'hc07c; // 0x20da
	13'h106e: q0 = 16'h000f; // 0x20dc
	13'h106f: q0 = 16'h48c0; // 0x20de
	13'h1070: q0 = 16'h2e00; // 0x20e0
	13'h1071: q0 = 16'h2007; // 0x20e2
	13'h1072: q0 = 16'h4281; // 0x20e4
	13'h1073: q0 = 16'h3205; // 0x20e6
	13'h1074: q0 = 16'he541; // 0x20e8
	13'h1075: q0 = 16'he3a0; // 0x20ea
	13'h1076: q0 = 16'h8194; // 0x20ec
	13'h1077: q0 = 16'h5245; // 0x20ee
	13'h1078: q0 = 16'h548d; // 0x20f0
	13'h1079: q0 = 16'h60de; // 0x20f2
	13'h107a: q0 = 16'h5246; // 0x20f4
	13'h107b: q0 = 16'h588c; // 0x20f6
	13'h107c: q0 = 16'h60c6; // 0x20f8
	13'h107d: q0 = 16'h4eb9; // 0x20fa
	13'h107e: q0 = 16'h0000; // 0x20fc
	13'h107f: q0 = 16'h2028; // 0x20fe
	13'h1080: q0 = 16'h3600; // 0x2100
	13'h1081: q0 = 16'h287c; // 0x2102
	13'h1082: q0 = 16'h0001; // 0x2104
	13'h1083: q0 = 16'h759a; // 0x2106
	13'h1084: q0 = 16'h4279; // 0x2108
	13'h1085: q0 = 16'h0001; // 0x210a
	13'h1086: q0 = 16'h7584; // 0x210c
	13'h1087: q0 = 16'h2a7c; // 0x210e
	13'h1088: q0 = 16'h0001; // 0x2110
	13'h1089: q0 = 16'h8684; // 0x2112
	13'h108a: q0 = 16'h4246; // 0x2114
	13'h108b: q0 = 16'hbc7c; // 0x2116
	13'h108c: q0 = 16'h000f; // 0x2118
	13'h108d: q0 = 16'h6c00; // 0x211a
	13'h108e: q0 = 16'h00b6; // 0x211c
	13'h108f: q0 = 16'h3006; // 0x211e
	13'h1090: q0 = 16'he540; // 0x2120
	13'h1091: q0 = 16'h48c0; // 0x2122
	13'h1092: q0 = 16'hd08b; // 0x2124
	13'h1093: q0 = 16'h2040; // 0x2126
	13'h1094: q0 = 16'h28a8; // 0x2128
	13'h1095: q0 = 16'h000a; // 0x212a
	13'h1096: q0 = 16'hbc7c; // 0x212c
	13'h1097: q0 = 16'h0003; // 0x212e
	13'h1098: q0 = 16'h6c38; // 0x2130
	13'h1099: q0 = 16'h3006; // 0x2132
	13'h109a: q0 = 16'he540; // 0x2134
	13'h109b: q0 = 16'h48c0; // 0x2136
	13'h109c: q0 = 16'hd08b; // 0x2138
	13'h109d: q0 = 16'h2040; // 0x213a
	13'h109e: q0 = 16'h3206; // 0x213c
	13'h109f: q0 = 16'he541; // 0x213e
	13'h10a0: q0 = 16'h48c1; // 0x2140
	13'h10a1: q0 = 16'hd2bc; // 0x2142
	13'h10a2: q0 = 16'h0001; // 0x2144
	13'h10a3: q0 = 16'h7f64; // 0x2146
	13'h10a4: q0 = 16'h2241; // 0x2148
	13'h10a5: q0 = 16'h22a8; // 0x214a
	13'h10a6: q0 = 16'h0046; // 0x214c
	13'h10a7: q0 = 16'h3006; // 0x214e
	13'h10a8: q0 = 16'he340; // 0x2150
	13'h10a9: q0 = 16'h48c0; // 0x2152
	13'h10aa: q0 = 16'hd0bc; // 0x2154
	13'h10ab: q0 = 16'h0001; // 0x2156
	13'h10ac: q0 = 16'h7efe; // 0x2158
	13'h10ad: q0 = 16'h2040; // 0x215a
	13'h10ae: q0 = 16'h3206; // 0x215c
	13'h10af: q0 = 16'he341; // 0x215e
	13'h10b0: q0 = 16'h48c1; // 0x2160
	13'h10b1: q0 = 16'hd28b; // 0x2162
	13'h10b2: q0 = 16'h2241; // 0x2164
	13'h10b3: q0 = 16'h30a9; // 0x2166
	13'h10b4: q0 = 16'h005c; // 0x2168
	13'h10b5: q0 = 16'hbc7c; // 0x216a
	13'h10b6: q0 = 16'h0009; // 0x216c
	13'h10b7: q0 = 16'h6c1a; // 0x216e
	13'h10b8: q0 = 16'h3006; // 0x2170
	13'h10b9: q0 = 16'h48c0; // 0x2172
	13'h10ba: q0 = 16'hd0bc; // 0x2174
	13'h10bb: q0 = 16'h0001; // 0x2176
	13'h10bc: q0 = 16'h7ba8; // 0x2178
	13'h10bd: q0 = 16'h2040; // 0x217a
	13'h10be: q0 = 16'h3406; // 0x217c
	13'h10bf: q0 = 16'h48c2; // 0x217e
	13'h10c0: q0 = 16'h220b; // 0x2180
	13'h10c1: q0 = 16'hd282; // 0x2182
	13'h10c2: q0 = 16'h2241; // 0x2184
	13'h10c3: q0 = 16'h10a9; // 0x2186
	13'h10c4: q0 = 16'h0052; // 0x2188
	13'h10c5: q0 = 16'hbc7c; // 0x218a
	13'h10c6: q0 = 16'h000a; // 0x218c
	13'h10c7: q0 = 16'h6c1c; // 0x218e
	13'h10c8: q0 = 16'h3006; // 0x2190
	13'h10c9: q0 = 16'he340; // 0x2192
	13'h10ca: q0 = 16'h48c0; // 0x2194
	13'h10cb: q0 = 16'hd0bc; // 0x2196
	13'h10cc: q0 = 16'h0001; // 0x2198
	13'h10cd: q0 = 16'h86b8; // 0x219a
	13'h10ce: q0 = 16'h2040; // 0x219c
	13'h10cf: q0 = 16'h3206; // 0x219e
	13'h10d0: q0 = 16'he341; // 0x21a0
	13'h10d1: q0 = 16'h48c1; // 0x21a2
	13'h10d2: q0 = 16'hd28b; // 0x21a4
	13'h10d3: q0 = 16'h2241; // 0x21a6
	13'h10d4: q0 = 16'h30a9; // 0x21a8
	13'h10d5: q0 = 16'h0062; // 0x21aa
	13'h10d6: q0 = 16'hbc7c; // 0x21ac
	13'h10d7: q0 = 16'h0008; // 0x21ae
	13'h10d8: q0 = 16'h6c16; // 0x21b0
	13'h10d9: q0 = 16'h3206; // 0x21b2
	13'h10da: q0 = 16'h48c1; // 0x21b4
	13'h10db: q0 = 16'h200b; // 0x21b6
	13'h10dc: q0 = 16'hd081; // 0x21b8
	13'h10dd: q0 = 16'h2040; // 0x21ba
	13'h10de: q0 = 16'h1028; // 0x21bc
	13'h10df: q0 = 16'h0076; // 0x21be
	13'h10e0: q0 = 16'h4880; // 0x21c0
	13'h10e1: q0 = 16'hc07c; // 0x21c2
	13'h10e2: q0 = 16'h00ff; // 0x21c4
	13'h10e3: q0 = 16'h3a80; // 0x21c6
	13'h10e4: q0 = 16'h5246; // 0x21c8
	13'h10e5: q0 = 16'h588c; // 0x21ca
	13'h10e6: q0 = 16'h548d; // 0x21cc
	13'h10e7: q0 = 16'h6000; // 0x21ce
	13'h10e8: q0 = 16'hff46; // 0x21d0
	13'h10e9: q0 = 16'h0803; // 0x21d2
	13'h10ea: q0 = 16'h0000; // 0x21d4
	13'h10eb: q0 = 16'h6706; // 0x21d6
	13'h10ec: q0 = 16'h4eb9; // 0x21d8
	13'h10ed: q0 = 16'h0000; // 0x21da
	13'h10ee: q0 = 16'haa34; // 0x21dc
	13'h10ef: q0 = 16'h0803; // 0x21de
	13'h10f0: q0 = 16'h0001; // 0x21e0
	13'h10f1: q0 = 16'h670c; // 0x21e2
	13'h10f2: q0 = 16'h42b9; // 0x21e4
	13'h10f3: q0 = 16'h0001; // 0x21e6
	13'h10f4: q0 = 16'h75ce; // 0x21e8
	13'h10f5: q0 = 16'h42b9; // 0x21ea
	13'h10f6: q0 = 16'h0001; // 0x21ec
	13'h10f7: q0 = 16'h75d2; // 0x21ee
	13'h10f8: q0 = 16'h0803; // 0x21f0
	13'h10f9: q0 = 16'h0002; // 0x21f2
	13'h10fa: q0 = 16'h6704; // 0x21f4
	13'h10fb: q0 = 16'h4245; // 0x21f6
	13'h10fc: q0 = 16'h6002; // 0x21f8
	13'h10fd: q0 = 16'h7a03; // 0x21fa
	13'h10fe: q0 = 16'h3e85; // 0x21fc
	13'h10ff: q0 = 16'h4eb9; // 0x21fe
	13'h1100: q0 = 16'h0000; // 0x2200
	13'h1101: q0 = 16'h55ce; // 0x2202
	13'h1102: q0 = 16'h0803; // 0x2204
	13'h1103: q0 = 16'h0003; // 0x2206
	13'h1104: q0 = 16'h6706; // 0x2208
	13'h1105: q0 = 16'h4eb9; // 0x220a
	13'h1106: q0 = 16'h0000; // 0x220c
	13'h1107: q0 = 16'h3cda; // 0x220e
	13'h1108: q0 = 16'h4eb9; // 0x2210
	13'h1109: q0 = 16'h0000; // 0x2212
	13'h110a: q0 = 16'hb2ae; // 0x2214
	13'h110b: q0 = 16'h0803; // 0x2216
	13'h110c: q0 = 16'h0004; // 0x2218
	13'h110d: q0 = 16'h671e; // 0x221a
	13'h110e: q0 = 16'h4246; // 0x221c
	13'h110f: q0 = 16'hbc7c; // 0x221e
	13'h1110: q0 = 16'h0008; // 0x2220
	13'h1111: q0 = 16'h6c16; // 0x2222
	13'h1112: q0 = 16'h3006; // 0x2224
	13'h1113: q0 = 16'he340; // 0x2226
	13'h1114: q0 = 16'h48c0; // 0x2228
	13'h1115: q0 = 16'hd0bc; // 0x222a
	13'h1116: q0 = 16'h0001; // 0x222c
	13'h1117: q0 = 16'h8684; // 0x222e
	13'h1118: q0 = 16'h2040; // 0x2230
	13'h1119: q0 = 16'h30bc; // 0x2232
	13'h111a: q0 = 16'h0080; // 0x2234
	13'h111b: q0 = 16'h5246; // 0x2236
	13'h111c: q0 = 16'h60e4; // 0x2238
	13'h111d: q0 = 16'h4a43; // 0x223a
	13'h111e: q0 = 16'h6704; // 0x223c
	13'h111f: q0 = 16'h4257; // 0x223e
	13'h1120: q0 = 16'h6004; // 0x2240
	13'h1121: q0 = 16'h3ebc; // 0x2242
	13'h1122: q0 = 16'h0001; // 0x2244
	13'h1123: q0 = 16'h0657; // 0x2246
	13'h1124: q0 = 16'h00b1; // 0x2248
	13'h1125: q0 = 16'h200e; // 0x224a
	13'h1126: q0 = 16'hd0bc; // 0x224c
	13'h1127: q0 = 16'hffff; // 0x224e
	13'h1128: q0 = 16'hffec; // 0x2250
	13'h1129: q0 = 16'h2f00; // 0x2252
	13'h112a: q0 = 16'h4eb9; // 0x2254
	13'h112b: q0 = 16'h0000; // 0x2256
	13'h112c: q0 = 16'h78f6; // 0x2258
	13'h112d: q0 = 16'h4a9f; // 0x225a
	13'h112e: q0 = 16'h4257; // 0x225c
	13'h112f: q0 = 16'h4267; // 0x225e
	13'h1130: q0 = 16'h3f3c; // 0x2260
	13'h1131: q0 = 16'h0001; // 0x2262
	13'h1132: q0 = 16'h3f3c; // 0x2264
	13'h1133: q0 = 16'h0011; // 0x2266
	13'h1134: q0 = 16'h200e; // 0x2268
	13'h1135: q0 = 16'hd0bc; // 0x226a
	13'h1136: q0 = 16'hffff; // 0x226c
	13'h1137: q0 = 16'hffec; // 0x226e
	13'h1138: q0 = 16'h2f00; // 0x2270
	13'h1139: q0 = 16'h4eb9; // 0x2272
	13'h113a: q0 = 16'h0000; // 0x2274
	13'h113b: q0 = 16'h026c; // 0x2276
	13'h113c: q0 = 16'hdefc; // 0x2278
	13'h113d: q0 = 16'h000a; // 0x227a
	13'h113e: q0 = 16'h4246; // 0x227c
	13'h113f: q0 = 16'h7a10; // 0x227e
	13'h1140: q0 = 16'hbc7c; // 0x2280
	13'h1141: q0 = 16'h0005; // 0x2282
	13'h1142: q0 = 16'h6c4a; // 0x2284
	13'h1143: q0 = 16'h3003; // 0x2286
	13'h1144: q0 = 16'h4281; // 0x2288
	13'h1145: q0 = 16'h3206; // 0x228a
	13'h1146: q0 = 16'he260; // 0x228c
	13'h1147: q0 = 16'hc07c; // 0x228e
	13'h1148: q0 = 16'h0001; // 0x2290
	13'h1149: q0 = 16'h6738; // 0x2292
	13'h114a: q0 = 16'h3e86; // 0x2294
	13'h114b: q0 = 16'h0657; // 0x2296
	13'h114c: q0 = 16'h00ac; // 0x2298
	13'h114d: q0 = 16'h200e; // 0x229a
	13'h114e: q0 = 16'hd0bc; // 0x229c
	13'h114f: q0 = 16'hffff; // 0x229e
	13'h1150: q0 = 16'hffec; // 0x22a0
	13'h1151: q0 = 16'h2f00; // 0x22a2
	13'h1152: q0 = 16'h4eb9; // 0x22a4
	13'h1153: q0 = 16'h0000; // 0x22a6
	13'h1154: q0 = 16'h78f6; // 0x22a8
	13'h1155: q0 = 16'h4a9f; // 0x22aa
	13'h1156: q0 = 16'h4257; // 0x22ac
	13'h1157: q0 = 16'h4267; // 0x22ae
	13'h1158: q0 = 16'h3f3c; // 0x22b0
	13'h1159: q0 = 16'h0004; // 0x22b2
	13'h115a: q0 = 16'h3f05; // 0x22b4
	13'h115b: q0 = 16'h5345; // 0x22b6
	13'h115c: q0 = 16'h200e; // 0x22b8
	13'h115d: q0 = 16'hd0bc; // 0x22ba
	13'h115e: q0 = 16'hffff; // 0x22bc
	13'h115f: q0 = 16'hffec; // 0x22be
	13'h1160: q0 = 16'h2f00; // 0x22c0
	13'h1161: q0 = 16'h4eb9; // 0x22c2
	13'h1162: q0 = 16'h0000; // 0x22c4
	13'h1163: q0 = 16'h026c; // 0x22c6
	13'h1164: q0 = 16'hdefc; // 0x22c8
	13'h1165: q0 = 16'h000a; // 0x22ca
	13'h1166: q0 = 16'h5246; // 0x22cc
	13'h1167: q0 = 16'h60b0; // 0x22ce
	13'h1168: q0 = 16'h4284; // 0x22d0
	13'h1169: q0 = 16'h2039; // 0x22d2
	13'h116a: q0 = 16'h0000; // 0x22d4
	13'h116b: q0 = 16'hc7d8; // 0x22d6
	13'h116c: q0 = 16'hb084; // 0x22d8
	13'h116d: q0 = 16'h6f1e; // 0x22da
	13'h116e: q0 = 16'h2a79; // 0x22dc
	13'h116f: q0 = 16'h0000; // 0x22de
	13'h1170: q0 = 16'hc7dc; // 0x22e0
	13'h1171: q0 = 16'h3c15; // 0x22e2
	13'h1172: q0 = 16'h2a79; // 0x22e4
	13'h1173: q0 = 16'h0000; // 0x22e6
	13'h1174: q0 = 16'hc7e0; // 0x22e8
	13'h1175: q0 = 16'h3c15; // 0x22ea
	13'h1176: q0 = 16'h0806; // 0x22ec
	13'h1177: q0 = 16'h0005; // 0x22ee
	13'h1178: q0 = 16'h6708; // 0x22f0
	13'h1179: q0 = 16'h4a43; // 0x22f2
	13'h117a: q0 = 16'h6602; // 0x22f4
	13'h117b: q0 = 16'h5284; // 0x22f6
	13'h117c: q0 = 16'h60d8; // 0x22f8
	13'h117d: q0 = 16'h4a9f; // 0x22fa
	13'h117e: q0 = 16'h4cdf; // 0x22fc
	13'h117f: q0 = 16'h38f8; // 0x22fe
	13'h1180: q0 = 16'h4e5e; // 0x2300
	13'h1181: q0 = 16'h4e75; // 0x2302
	13'h1182: q0 = 16'h4e56; // 0x2304
	13'h1183: q0 = 16'h0000; // 0x2306
	13'h1184: q0 = 16'h48e7; // 0x2308
	13'h1185: q0 = 16'h071c; // 0x230a
	13'h1186: q0 = 16'h267c; // 0x230c
	13'h1187: q0 = 16'h0001; // 0x230e
	13'h1188: q0 = 16'h7fd4; // 0x2310
	13'h1189: q0 = 16'h4eb9; // 0x2312
	13'h118a: q0 = 16'h0000; // 0x2314
	13'h118b: q0 = 16'h1564; // 0x2316
	13'h118c: q0 = 16'h287c; // 0x2318
	13'h118d: q0 = 16'h0001; // 0x231a
	13'h118e: q0 = 16'h759a; // 0x231c
	13'h118f: q0 = 16'h2a7c; // 0x231e
	13'h1190: q0 = 16'h0001; // 0x2320
	13'h1191: q0 = 16'h8684; // 0x2322
	13'h1192: q0 = 16'h4247; // 0x2324
	13'h1193: q0 = 16'hbe7c; // 0x2326
	13'h1194: q0 = 16'h000f; // 0x2328
	13'h1195: q0 = 16'h6c00; // 0x232a
	13'h1196: q0 = 16'h00b0; // 0x232c
	13'h1197: q0 = 16'h3007; // 0x232e
	13'h1198: q0 = 16'he540; // 0x2330
	13'h1199: q0 = 16'h48c0; // 0x2332
	13'h119a: q0 = 16'hd08b; // 0x2334
	13'h119b: q0 = 16'h2040; // 0x2336
	13'h119c: q0 = 16'h2154; // 0x2338
	13'h119d: q0 = 16'h000a; // 0x233a
	13'h119e: q0 = 16'hbe7c; // 0x233c
	13'h119f: q0 = 16'h0003; // 0x233e
	13'h11a0: q0 = 16'h6c38; // 0x2340
	13'h11a1: q0 = 16'h3007; // 0x2342
	13'h11a2: q0 = 16'he540; // 0x2344
	13'h11a3: q0 = 16'h48c0; // 0x2346
	13'h11a4: q0 = 16'hd0bc; // 0x2348
	13'h11a5: q0 = 16'h0001; // 0x234a
	13'h11a6: q0 = 16'h7f64; // 0x234c
	13'h11a7: q0 = 16'h2040; // 0x234e
	13'h11a8: q0 = 16'h3207; // 0x2350
	13'h11a9: q0 = 16'he541; // 0x2352
	13'h11aa: q0 = 16'h48c1; // 0x2354
	13'h11ab: q0 = 16'hd28b; // 0x2356
	13'h11ac: q0 = 16'h2241; // 0x2358
	13'h11ad: q0 = 16'h2350; // 0x235a
	13'h11ae: q0 = 16'h0046; // 0x235c
	13'h11af: q0 = 16'h3007; // 0x235e
	13'h11b0: q0 = 16'he340; // 0x2360
	13'h11b1: q0 = 16'h48c0; // 0x2362
	13'h11b2: q0 = 16'hd08b; // 0x2364
	13'h11b3: q0 = 16'h2040; // 0x2366
	13'h11b4: q0 = 16'h3207; // 0x2368
	13'h11b5: q0 = 16'he341; // 0x236a
	13'h11b6: q0 = 16'h48c1; // 0x236c
	13'h11b7: q0 = 16'hd2bc; // 0x236e
	13'h11b8: q0 = 16'h0001; // 0x2370
	13'h11b9: q0 = 16'h7efe; // 0x2372
	13'h11ba: q0 = 16'h2241; // 0x2374
	13'h11bb: q0 = 16'h3151; // 0x2376
	13'h11bc: q0 = 16'h005c; // 0x2378
	13'h11bd: q0 = 16'hbe7c; // 0x237a
	13'h11be: q0 = 16'h0009; // 0x237c
	13'h11bf: q0 = 16'h6c1a; // 0x237e
	13'h11c0: q0 = 16'h3207; // 0x2380
	13'h11c1: q0 = 16'h48c1; // 0x2382
	13'h11c2: q0 = 16'h200b; // 0x2384
	13'h11c3: q0 = 16'hd081; // 0x2386
	13'h11c4: q0 = 16'h2040; // 0x2388
	13'h11c5: q0 = 16'h3207; // 0x238a
	13'h11c6: q0 = 16'h48c1; // 0x238c
	13'h11c7: q0 = 16'hd2bc; // 0x238e
	13'h11c8: q0 = 16'h0001; // 0x2390
	13'h11c9: q0 = 16'h7ba8; // 0x2392
	13'h11ca: q0 = 16'h2241; // 0x2394
	13'h11cb: q0 = 16'h1151; // 0x2396
	13'h11cc: q0 = 16'h0052; // 0x2398
	13'h11cd: q0 = 16'hbe7c; // 0x239a
	13'h11ce: q0 = 16'h000a; // 0x239c
	13'h11cf: q0 = 16'h6c1c; // 0x239e
	13'h11d0: q0 = 16'h3007; // 0x23a0
	13'h11d1: q0 = 16'he340; // 0x23a2
	13'h11d2: q0 = 16'h48c0; // 0x23a4
	13'h11d3: q0 = 16'hd08b; // 0x23a6
	13'h11d4: q0 = 16'h2040; // 0x23a8
	13'h11d5: q0 = 16'h3207; // 0x23aa
	13'h11d6: q0 = 16'he341; // 0x23ac
	13'h11d7: q0 = 16'h48c1; // 0x23ae
	13'h11d8: q0 = 16'hd2bc; // 0x23b0
	13'h11d9: q0 = 16'h0001; // 0x23b2
	13'h11da: q0 = 16'h86b8; // 0x23b4
	13'h11db: q0 = 16'h2241; // 0x23b6
	13'h11dc: q0 = 16'h3151; // 0x23b8
	13'h11dd: q0 = 16'h0062; // 0x23ba
	13'h11de: q0 = 16'hbe7c; // 0x23bc
	13'h11df: q0 = 16'h0008; // 0x23be
	13'h11e0: q0 = 16'h6c10; // 0x23c0
	13'h11e1: q0 = 16'h3207; // 0x23c2
	13'h11e2: q0 = 16'h48c1; // 0x23c4
	13'h11e3: q0 = 16'h200b; // 0x23c6
	13'h11e4: q0 = 16'hd081; // 0x23c8
	13'h11e5: q0 = 16'h2040; // 0x23ca
	13'h11e6: q0 = 16'h3215; // 0x23cc
	13'h11e7: q0 = 16'h1141; // 0x23ce
	13'h11e8: q0 = 16'h0076; // 0x23d0
	13'h11e9: q0 = 16'h5247; // 0x23d2
	13'h11ea: q0 = 16'h588c; // 0x23d4
	13'h11eb: q0 = 16'h548d; // 0x23d6
	13'h11ec: q0 = 16'h6000; // 0x23d8
	13'h11ed: q0 = 16'hff4c; // 0x23da
	13'h11ee: q0 = 16'h4eb9; // 0x23dc
	13'h11ef: q0 = 16'h0000; // 0x23de
	13'h11f0: q0 = 16'h2028; // 0x23e0
	13'h11f1: q0 = 16'h287c; // 0x23e2
	13'h11f2: q0 = 16'h0001; // 0x23e4
	13'h11f3: q0 = 16'h7fd4; // 0x23e6
	13'h11f4: q0 = 16'h2a79; // 0x23e8
	13'h11f5: q0 = 16'h0000; // 0x23ea
	13'h11f6: q0 = 16'hc7e4; // 0x23ec
	13'h11f7: q0 = 16'h4247; // 0x23ee
	13'h11f8: q0 = 16'hbe7c; // 0x23f0
	13'h11f9: q0 = 16'h0020; // 0x23f2
	13'h11fa: q0 = 16'h6c30; // 0x23f4
	13'h11fb: q0 = 16'h2014; // 0x23f6
	13'h11fc: q0 = 16'hc0bc; // 0x23f8
	13'h11fd: q0 = 16'h0000; // 0x23fa
	13'h11fe: q0 = 16'h000f; // 0x23fc
	13'h11ff: q0 = 16'h3ac0; // 0x23fe
	13'h1200: q0 = 16'h7c01; // 0x2400
	13'h1201: q0 = 16'hbc7c; // 0x2402
	13'h1202: q0 = 16'h0008; // 0x2404
	13'h1203: q0 = 16'h6c18; // 0x2406
	13'h1204: q0 = 16'h2014; // 0x2408
	13'h1205: q0 = 16'h4281; // 0x240a
	13'h1206: q0 = 16'h3206; // 0x240c
	13'h1207: q0 = 16'he541; // 0x240e
	13'h1208: q0 = 16'he2a0; // 0x2410
	13'h1209: q0 = 16'hc0bc; // 0x2412
	13'h120a: q0 = 16'h0000; // 0x2414
	13'h120b: q0 = 16'h000f; // 0x2416
	13'h120c: q0 = 16'h3a80; // 0x2418
	13'h120d: q0 = 16'h5246; // 0x241a
	13'h120e: q0 = 16'h548d; // 0x241c
	13'h120f: q0 = 16'h60e2; // 0x241e
	13'h1210: q0 = 16'h5247; // 0x2420
	13'h1211: q0 = 16'h588c; // 0x2422
	13'h1212: q0 = 16'h60ca; // 0x2424
	13'h1213: q0 = 16'h0079; // 0x2426
	13'h1214: q0 = 16'h0002; // 0x2428
	13'h1215: q0 = 16'h0001; // 0x242a
	13'h1216: q0 = 16'h861e; // 0x242c
	13'h1217: q0 = 16'h4a9f; // 0x242e
	13'h1218: q0 = 16'h4cdf; // 0x2430
	13'h1219: q0 = 16'h38c0; // 0x2432
	13'h121a: q0 = 16'h4e5e; // 0x2434
	13'h121b: q0 = 16'h4e75; // 0x2436
	13'h121c: q0 = 16'h4e56; // 0x2438
	13'h121d: q0 = 16'hffe8; // 0x243a
	13'h121e: q0 = 16'h48e7; // 0x243c
	13'h121f: q0 = 16'h0304; // 0x243e
	13'h1220: q0 = 16'h2a6e; // 0x2440
	13'h1221: q0 = 16'h0008; // 0x2442
	13'h1222: q0 = 16'h4eb9; // 0x2444
	13'h1223: q0 = 16'h0000; // 0x2446
	13'h1224: q0 = 16'h4ec6; // 0x2448
	13'h1225: q0 = 16'hb07c; // 0x244a
	13'h1226: q0 = 16'h0005; // 0x244c
	13'h1227: q0 = 16'h6674; // 0x244e
	13'h1228: q0 = 16'h082d; // 0x2450
	13'h1229: q0 = 16'h0005; // 0x2452
	13'h122a: q0 = 16'h000f; // 0x2454
	13'h122b: q0 = 16'h666c; // 0x2456
	13'h122c: q0 = 16'h006d; // 0x2458
	13'h122d: q0 = 16'h0020; // 0x245a
	13'h122e: q0 = 16'h000e; // 0x245c
	13'h122f: q0 = 16'h206d; // 0x245e
	13'h1230: q0 = 16'h001e; // 0x2460
	13'h1231: q0 = 16'h3ea8; // 0x2462
	13'h1232: q0 = 16'h0002; // 0x2464
	13'h1233: q0 = 16'h4eb9; // 0x2466
	13'h1234: q0 = 16'h0000; // 0x2468
	13'h1235: q0 = 16'h4f30; // 0x246a
	13'h1236: q0 = 16'h9157; // 0x246c
	13'h1237: q0 = 16'h206d; // 0x246e
	13'h1238: q0 = 16'h001e; // 0x2470
	13'h1239: q0 = 16'h3f10; // 0x2472
	13'h123a: q0 = 16'h4eb9; // 0x2474
	13'h123b: q0 = 16'h0000; // 0x2476
	13'h123c: q0 = 16'h4ee2; // 0x2478
	13'h123d: q0 = 16'h9157; // 0x247a
	13'h123e: q0 = 16'h4eb9; // 0x247c
	13'h123f: q0 = 16'h0000; // 0x247e
	13'h1240: q0 = 16'h0a1c; // 0x2480
	13'h1241: q0 = 16'h4a5f; // 0x2482
	13'h1242: q0 = 16'h3a80; // 0x2484
	13'h1243: q0 = 16'h302d; // 0x2486
	13'h1244: q0 = 16'h000e; // 0x2488
	13'h1245: q0 = 16'hc07c; // 0x248a
	13'h1246: q0 = 16'h000f; // 0x248c
	13'h1247: q0 = 16'hb07c; // 0x248e
	13'h1248: q0 = 16'h0001; // 0x2490
	13'h1249: q0 = 16'h6708; // 0x2492
	13'h124a: q0 = 16'he0ed; // 0x2494
	13'h124b: q0 = 16'h000c; // 0x2496
	13'h124c: q0 = 16'h426d; // 0x2498
	13'h124d: q0 = 16'h000a; // 0x249a
	13'h124e: q0 = 16'he1ed; // 0x249c
	13'h124f: q0 = 16'h0002; // 0x249e
	13'h1250: q0 = 16'h3ead; // 0x24a0
	13'h1251: q0 = 16'h0002; // 0x24a2
	13'h1252: q0 = 16'h3f15; // 0x24a4
	13'h1253: q0 = 16'h4eb9; // 0x24a6
	13'h1254: q0 = 16'h0000; // 0x24a8
	13'h1255: q0 = 16'h1280; // 0x24aa
	13'h1256: q0 = 16'h4a5f; // 0x24ac
	13'h1257: q0 = 16'h3b40; // 0x24ae
	13'h1258: q0 = 16'h0004; // 0x24b0
	13'h1259: q0 = 16'h3ead; // 0x24b2
	13'h125a: q0 = 16'h0002; // 0x24b4
	13'h125b: q0 = 16'h3f15; // 0x24b6
	13'h125c: q0 = 16'h4eb9; // 0x24b8
	13'h125d: q0 = 16'h0000; // 0x24ba
	13'h125e: q0 = 16'ha730; // 0x24bc
	13'h125f: q0 = 16'h4a5f; // 0x24be
	13'h1260: q0 = 16'h3b40; // 0x24c0
	13'h1261: q0 = 16'h0006; // 0x24c2
	13'h1262: q0 = 16'h302d; // 0x24c4
	13'h1263: q0 = 16'h000e; // 0x24c6
	13'h1264: q0 = 16'hc07c; // 0x24c8
	13'h1265: q0 = 16'h000f; // 0x24ca
	13'h1266: q0 = 16'hb07c; // 0x24cc
	13'h1267: q0 = 16'h0001; // 0x24ce
	13'h1268: q0 = 16'h6700; // 0x24d0
	13'h1269: q0 = 16'h043e; // 0x24d2
	13'h126a: q0 = 16'h4a79; // 0x24d4
	13'h126b: q0 = 16'h0001; // 0x24d6
	13'h126c: q0 = 16'h75e6; // 0x24d8
	13'h126d: q0 = 16'h673c; // 0x24da
	13'h126e: q0 = 16'h2d79; // 0x24dc
	13'h126f: q0 = 16'h0000; // 0x24de
	13'h1270: q0 = 16'hc80c; // 0x24e0
	13'h1271: q0 = 16'hffe8; // 0x24e2
	13'h1272: q0 = 16'h06ae; // 0x24e4
	13'h1273: q0 = 16'h0000; // 0x24e6
	13'h1274: q0 = 16'h7000; // 0x24e8
	13'h1275: q0 = 16'hffe8; // 0x24ea
	13'h1276: q0 = 16'h206e; // 0x24ec
	13'h1277: q0 = 16'hffe8; // 0x24ee
	13'h1278: q0 = 16'h2010; // 0x24f0
	13'h1279: q0 = 16'hc0bc; // 0x24f2
	13'h127a: q0 = 16'h0000; // 0x24f4
	13'h127b: q0 = 16'h003f; // 0x24f6
	13'h127c: q0 = 16'h661e; // 0x24f8
	13'h127d: q0 = 16'h206e; // 0x24fa
	13'h127e: q0 = 16'hffe8; // 0x24fc
	13'h127f: q0 = 16'h4a90; // 0x24fe
	13'h1280: q0 = 16'h6f16; // 0x2500
	13'h1281: q0 = 16'h206e; // 0x2502
	13'h1282: q0 = 16'hffe8; // 0x2504
	13'h1283: q0 = 16'h5290; // 0x2506
	13'h1284: q0 = 16'h2d6e; // 0x2508
	13'h1285: q0 = 16'hffe8; // 0x250a
	13'h1286: q0 = 16'hffec; // 0x250c
	13'h1287: q0 = 16'h206e; // 0x250e
	13'h1288: q0 = 16'hffec; // 0x2510
	13'h1289: q0 = 16'h317c; // 0x2512
	13'h128a: q0 = 16'h0001; // 0x2514
	13'h128b: q0 = 16'hffd6; // 0x2516
	13'h128c: q0 = 16'h4a6d; // 0x2518
	13'h128d: q0 = 16'h0014; // 0x251a
	13'h128e: q0 = 16'h6f04; // 0x251c
	13'h128f: q0 = 16'h536d; // 0x251e
	13'h1290: q0 = 16'h0014; // 0x2520
	13'h1291: q0 = 16'h4a6d; // 0x2522
	13'h1292: q0 = 16'h0014; // 0x2524
	13'h1293: q0 = 16'h6600; // 0x2526
	13'h1294: q0 = 16'h00ca; // 0x2528
	13'h1295: q0 = 16'h082d; // 0x252a
	13'h1296: q0 = 16'h0004; // 0x252c
	13'h1297: q0 = 16'h000f; // 0x252e
	13'h1298: q0 = 16'h6600; // 0x2530
	13'h1299: q0 = 16'h00c0; // 0x2532
	13'h129a: q0 = 16'h206d; // 0x2534
	13'h129b: q0 = 16'h001e; // 0x2536
	13'h129c: q0 = 16'h3d50; // 0x2538
	13'h129d: q0 = 16'hfffe; // 0x253a
	13'h129e: q0 = 16'h206d; // 0x253c
	13'h129f: q0 = 16'h001e; // 0x253e
	13'h12a0: q0 = 16'h3d68; // 0x2540
	13'h12a1: q0 = 16'h0002; // 0x2542
	13'h12a2: q0 = 16'hfffc; // 0x2544
	13'h12a3: q0 = 16'h4257; // 0x2546
	13'h12a4: q0 = 16'h200e; // 0x2548
	13'h12a5: q0 = 16'hd0bc; // 0x254a
	13'h12a6: q0 = 16'hffff; // 0x254c
	13'h12a7: q0 = 16'hfffc; // 0x254e
	13'h12a8: q0 = 16'h2f00; // 0x2550
	13'h12a9: q0 = 16'h200e; // 0x2552
	13'h12aa: q0 = 16'hd0bc; // 0x2554
	13'h12ab: q0 = 16'hffff; // 0x2556
	13'h12ac: q0 = 16'hfffe; // 0x2558
	13'h12ad: q0 = 16'h2f00; // 0x255a
	13'h12ae: q0 = 16'h4eb9; // 0x255c
	13'h12af: q0 = 16'h0000; // 0x255e
	13'h12b0: q0 = 16'h5d44; // 0x2560
	13'h12b1: q0 = 16'hbf8f; // 0x2562
	13'h12b2: q0 = 16'h4a40; // 0x2564
	13'h12b3: q0 = 16'h6700; // 0x2566
	13'h12b4: q0 = 16'h008a; // 0x2568
	13'h12b5: q0 = 16'h3ebc; // 0x256a
	13'h12b6: q0 = 16'h0002; // 0x256c
	13'h12b7: q0 = 16'h4eb9; // 0x256e
	13'h12b8: q0 = 16'h0000; // 0x2570
	13'h12b9: q0 = 16'h8ee8; // 0x2572
	13'h12ba: q0 = 16'h4a79; // 0x2574
	13'h12bb: q0 = 16'h0001; // 0x2576
	13'h12bc: q0 = 16'h8676; // 0x2578
	13'h12bd: q0 = 16'h661c; // 0x257a
	13'h12be: q0 = 16'h206d; // 0x257c
	13'h12bf: q0 = 16'h001a; // 0x257e
	13'h12c0: q0 = 16'h3010; // 0x2580
	13'h12c1: q0 = 16'h5340; // 0x2582
	13'h12c2: q0 = 16'he540; // 0x2584
	13'h12c3: q0 = 16'h48c0; // 0x2586
	13'h12c4: q0 = 16'hd0bc; // 0x2588
	13'h12c5: q0 = 16'h0000; // 0x258a
	13'h12c6: q0 = 16'hc7e8; // 0x258c
	13'h12c7: q0 = 16'h2040; // 0x258e
	13'h12c8: q0 = 16'h2e90; // 0x2590
	13'h12c9: q0 = 16'h4eb9; // 0x2592
	13'h12ca: q0 = 16'h0000; // 0x2594
	13'h12cb: q0 = 16'h7dd8; // 0x2596
	13'h12cc: q0 = 16'h3eae; // 0x2598
	13'h12cd: q0 = 16'hfffc; // 0x259a
	13'h12ce: q0 = 16'h3f2e; // 0x259c
	13'h12cf: q0 = 16'hfffe; // 0x259e
	13'h12d0: q0 = 16'h2f0d; // 0x25a0
	13'h12d1: q0 = 16'h4eb9; // 0x25a2
	13'h12d2: q0 = 16'h0000; // 0x25a4
	13'h12d3: q0 = 16'h2dc2; // 0x25a6
	13'h12d4: q0 = 16'h5c4f; // 0x25a8
	13'h12d5: q0 = 16'h3b6e; // 0x25aa
	13'h12d6: q0 = 16'hfffc; // 0x25ac
	13'h12d7: q0 = 16'h0018; // 0x25ae
	13'h12d8: q0 = 16'h206d; // 0x25b0
	13'h12d9: q0 = 16'h001e; // 0x25b2
	13'h12da: q0 = 16'h317c; // 0x25b4
	13'h12db: q0 = 16'h0017; // 0x25b6
	13'h12dc: q0 = 16'h0006; // 0x25b8
	13'h12dd: q0 = 16'h206d; // 0x25ba
	13'h12de: q0 = 16'h0026; // 0x25bc
	13'h12df: q0 = 16'h317c; // 0x25be
	13'h12e0: q0 = 16'h0017; // 0x25c0
	13'h12e1: q0 = 16'h0006; // 0x25c2
	13'h12e2: q0 = 16'h3b7c; // 0x25c4
	13'h12e3: q0 = 16'h0001; // 0x25c6
	13'h12e4: q0 = 16'h0008; // 0x25c8
	13'h12e5: q0 = 16'h4aad; // 0x25ca
	13'h12e6: q0 = 16'h0010; // 0x25cc
	13'h12e7: q0 = 16'h670e; // 0x25ce
	13'h12e8: q0 = 16'h2ead; // 0x25d0
	13'h12e9: q0 = 16'h0010; // 0x25d2
	13'h12ea: q0 = 16'h4eb9; // 0x25d4
	13'h12eb: q0 = 16'h0000; // 0x25d6
	13'h12ec: q0 = 16'h3356; // 0x25d8
	13'h12ed: q0 = 16'h42ad; // 0x25da
	13'h12ee: q0 = 16'h0010; // 0x25dc
	13'h12ef: q0 = 16'h302d; // 0x25de
	13'h12f0: q0 = 16'h000e; // 0x25e0
	13'h12f1: q0 = 16'hc07c; // 0x25e2
	13'h12f2: q0 = 16'hf000; // 0x25e4
	13'h12f3: q0 = 16'h807c; // 0x25e6
	13'h12f4: q0 = 16'h0003; // 0x25e8
	13'h12f5: q0 = 16'h3b40; // 0x25ea
	13'h12f6: q0 = 16'h000e; // 0x25ec
	13'h12f7: q0 = 16'h6000; // 0x25ee
	13'h12f8: q0 = 16'h0320; // 0x25f0
	13'h12f9: q0 = 16'h200e; // 0x25f2
	13'h12fa: q0 = 16'hd0bc; // 0x25f4
	13'h12fb: q0 = 16'hffff; // 0x25f6
	13'h12fc: q0 = 16'hfff0; // 0x25f8
	13'h12fd: q0 = 16'h2e80; // 0x25fa
	13'h12fe: q0 = 16'h200e; // 0x25fc
	13'h12ff: q0 = 16'hd0bc; // 0x25fe
	13'h1300: q0 = 16'hffff; // 0x2600
	13'h1301: q0 = 16'hfff2; // 0x2602
	13'h1302: q0 = 16'h2f00; // 0x2604
	13'h1303: q0 = 16'h200e; // 0x2606
	13'h1304: q0 = 16'hd0bc; // 0x2608
	13'h1305: q0 = 16'hffff; // 0x260a
	13'h1306: q0 = 16'hfff4; // 0x260c
	13'h1307: q0 = 16'h2f00; // 0x260e
	13'h1308: q0 = 16'h200e; // 0x2610
	13'h1309: q0 = 16'hd0bc; // 0x2612
	13'h130a: q0 = 16'hffff; // 0x2614
	13'h130b: q0 = 16'hfff6; // 0x2616
	13'h130c: q0 = 16'h2f00; // 0x2618
	13'h130d: q0 = 16'h2f0d; // 0x261a
	13'h130e: q0 = 16'h206d; // 0x261c
	13'h130f: q0 = 16'h001e; // 0x261e
	13'h1310: q0 = 16'h3f28; // 0x2620
	13'h1311: q0 = 16'h0002; // 0x2622
	13'h1312: q0 = 16'h206d; // 0x2624
	13'h1313: q0 = 16'h001e; // 0x2626
	13'h1314: q0 = 16'h3f10; // 0x2628
	13'h1315: q0 = 16'h4eb9; // 0x262a
	13'h1316: q0 = 16'h0000; // 0x262c
	13'h1317: q0 = 16'h36d8; // 0x262e
	13'h1318: q0 = 16'hdefc; // 0x2630
	13'h1319: q0 = 16'h0014; // 0x2632
	13'h131a: q0 = 16'h2d40; // 0x2634
	13'h131b: q0 = 16'hfff8; // 0x2636
	13'h131c: q0 = 16'h4aae; // 0x2638
	13'h131d: q0 = 16'hfff8; // 0x263a
	13'h131e: q0 = 16'h665e; // 0x263c
	13'h131f: q0 = 16'h206d; // 0x263e
	13'h1320: q0 = 16'h001a; // 0x2640
	13'h1321: q0 = 16'h0c50; // 0x2642
	13'h1322: q0 = 16'h0002; // 0x2644
	13'h1323: q0 = 16'h670a; // 0x2646
	13'h1324: q0 = 16'h206d; // 0x2648
	13'h1325: q0 = 16'h001a; // 0x264a
	13'h1326: q0 = 16'h0c50; // 0x264c
	13'h1327: q0 = 16'h0003; // 0x264e
	13'h1328: q0 = 16'h664a; // 0x2650
	13'h1329: q0 = 16'h200e; // 0x2652
	13'h132a: q0 = 16'hd0bc; // 0x2654
	13'h132b: q0 = 16'hffff; // 0x2656
	13'h132c: q0 = 16'hfff0; // 0x2658
	13'h132d: q0 = 16'h2e80; // 0x265a
	13'h132e: q0 = 16'h200e; // 0x265c
	13'h132f: q0 = 16'hd0bc; // 0x265e
	13'h1330: q0 = 16'hffff; // 0x2660
	13'h1331: q0 = 16'hfff2; // 0x2662
	13'h1332: q0 = 16'h2f00; // 0x2664
	13'h1333: q0 = 16'h200e; // 0x2666
	13'h1334: q0 = 16'hd0bc; // 0x2668
	13'h1335: q0 = 16'hffff; // 0x266a
	13'h1336: q0 = 16'hfff4; // 0x266c
	13'h1337: q0 = 16'h2f00; // 0x266e
	13'h1338: q0 = 16'h200e; // 0x2670
	13'h1339: q0 = 16'hd0bc; // 0x2672
	13'h133a: q0 = 16'hffff; // 0x2674
	13'h133b: q0 = 16'hfff6; // 0x2676
	13'h133c: q0 = 16'h2f00; // 0x2678
	13'h133d: q0 = 16'h2f0d; // 0x267a
	13'h133e: q0 = 16'h206d; // 0x267c
	13'h133f: q0 = 16'h001e; // 0x267e
	13'h1340: q0 = 16'h3f28; // 0x2680
	13'h1341: q0 = 16'h0002; // 0x2682
	13'h1342: q0 = 16'h0657; // 0x2684
	13'h1343: q0 = 16'h0200; // 0x2686
	13'h1344: q0 = 16'h206d; // 0x2688
	13'h1345: q0 = 16'h001e; // 0x268a
	13'h1346: q0 = 16'h3f10; // 0x268c
	13'h1347: q0 = 16'h4eb9; // 0x268e
	13'h1348: q0 = 16'h0000; // 0x2690
	13'h1349: q0 = 16'h36d8; // 0x2692
	13'h134a: q0 = 16'hdefc; // 0x2694
	13'h134b: q0 = 16'h0014; // 0x2696
	13'h134c: q0 = 16'h2d40; // 0x2698
	13'h134d: q0 = 16'hfff8; // 0x269a
	13'h134e: q0 = 16'h4aae; // 0x269c
	13'h134f: q0 = 16'hfff8; // 0x269e
	13'h1350: q0 = 16'h6700; // 0x26a0
	13'h1351: q0 = 16'h026a; // 0x26a2
	13'h1352: q0 = 16'h4aad; // 0x26a4
	13'h1353: q0 = 16'h0010; // 0x26a6
	13'h1354: q0 = 16'h670e; // 0x26a8
	13'h1355: q0 = 16'h2ead; // 0x26aa
	13'h1356: q0 = 16'h0010; // 0x26ac
	13'h1357: q0 = 16'h4eb9; // 0x26ae
	13'h1358: q0 = 16'h0000; // 0x26b0
	13'h1359: q0 = 16'h3356; // 0x26b2
	13'h135a: q0 = 16'h42ad; // 0x26b4
	13'h135b: q0 = 16'h0010; // 0x26b6
	13'h135c: q0 = 16'h082d; // 0x26b8
	13'h135d: q0 = 16'h0004; // 0x26ba
	13'h135e: q0 = 16'h000f; // 0x26bc
	13'h135f: q0 = 16'h6630; // 0x26be
	13'h1360: q0 = 16'h082d; // 0x26c0
	13'h1361: q0 = 16'h0005; // 0x26c2
	13'h1362: q0 = 16'h000f; // 0x26c4
	13'h1363: q0 = 16'h6628; // 0x26c6
	13'h1364: q0 = 16'h3aae; // 0x26c8
	13'h1365: q0 = 16'hfff4; // 0x26ca
	13'h1366: q0 = 16'h3b6e; // 0x26cc
	13'h1367: q0 = 16'hfff2; // 0x26ce
	13'h1368: q0 = 16'h0004; // 0x26d0
	13'h1369: q0 = 16'h3b6e; // 0x26d2
	13'h136a: q0 = 16'hfff0; // 0x26d4
	13'h136b: q0 = 16'h0006; // 0x26d6
	13'h136c: q0 = 16'h0c6d; // 0x26d8
	13'h136d: q0 = 16'h0001; // 0x26da
	13'h136e: q0 = 16'h000c; // 0x26dc
	13'h136f: q0 = 16'h6e06; // 0x26de
	13'h1370: q0 = 16'h426d; // 0x26e0
	13'h1371: q0 = 16'h000c; // 0x26e2
	13'h1372: q0 = 16'h6006; // 0x26e4
	13'h1373: q0 = 16'h3b7c; // 0x26e6
	13'h1374: q0 = 16'h0001; // 0x26e8
	13'h1375: q0 = 16'h000c; // 0x26ea
	13'h1376: q0 = 16'h426d; // 0x26ec
	13'h1377: q0 = 16'h000a; // 0x26ee
	13'h1378: q0 = 16'h082d; // 0x26f0
	13'h1379: q0 = 16'h0004; // 0x26f2
	13'h137a: q0 = 16'h000f; // 0x26f4
	13'h137b: q0 = 16'h6704; // 0x26f6
	13'h137c: q0 = 16'h7e03; // 0x26f8
	13'h137d: q0 = 16'h6016; // 0x26fa
	13'h137e: q0 = 16'h3039; // 0x26fc
	13'h137f: q0 = 16'h0001; // 0x26fe
	13'h1380: q0 = 16'h8a76; // 0x2700
	13'h1381: q0 = 16'h226d; // 0x2702
	13'h1382: q0 = 16'h001a; // 0x2704
	13'h1383: q0 = 16'h4281; // 0x2706
	13'h1384: q0 = 16'h3211; // 0x2708
	13'h1385: q0 = 16'he260; // 0x270a
	13'h1386: q0 = 16'h3e00; // 0x270c
	13'h1387: q0 = 16'hce7c; // 0x270e
	13'h1388: q0 = 16'h0007; // 0x2710
	13'h1389: q0 = 16'h3007; // 0x2712
	13'h138a: q0 = 16'h6000; // 0x2714
	13'h138b: q0 = 16'h00da; // 0x2716
	13'h138c: q0 = 16'h302d; // 0x2718
	13'h138d: q0 = 16'h000e; // 0x271a
	13'h138e: q0 = 16'h807c; // 0x271c
	13'h138f: q0 = 16'h0100; // 0x271e
	13'h1390: q0 = 16'h3b40; // 0x2720
	13'h1391: q0 = 16'h000e; // 0x2722
	13'h1392: q0 = 16'h6000; // 0x2724
	13'h1393: q0 = 16'h00de; // 0x2726
	13'h1394: q0 = 16'h206d; // 0x2728
	13'h1395: q0 = 16'h0022; // 0x272a
	13'h1396: q0 = 16'h317c; // 0x272c
	13'h1397: q0 = 16'h0059; // 0x272e
	13'h1398: q0 = 16'h0004; // 0x2730
	13'h1399: q0 = 16'h6000; // 0x2732
	13'h139a: q0 = 16'h00d0; // 0x2734
	13'h139b: q0 = 16'h206d; // 0x2736
	13'h139c: q0 = 16'h0022; // 0x2738
	13'h139d: q0 = 16'h317c; // 0x273a
	13'h139e: q0 = 16'h0058; // 0x273c
	13'h139f: q0 = 16'h0004; // 0x273e
	13'h13a0: q0 = 16'h206d; // 0x2740
	13'h13a1: q0 = 16'h0022; // 0x2742
	13'h13a2: q0 = 16'h317c; // 0x2744
	13'h13a3: q0 = 16'h0010; // 0x2746
	13'h13a4: q0 = 16'h0006; // 0x2748
	13'h13a5: q0 = 16'h6000; // 0x274a
	13'h13a6: q0 = 16'h00b8; // 0x274c
	13'h13a7: q0 = 16'h302d; // 0x274e
	13'h13a8: q0 = 16'h000e; // 0x2750
	13'h13a9: q0 = 16'h807c; // 0x2752
	13'h13aa: q0 = 16'h0400; // 0x2754
	13'h13ab: q0 = 16'h3b40; // 0x2756
	13'h13ac: q0 = 16'h000e; // 0x2758
	13'h13ad: q0 = 16'h6000; // 0x275a
	13'h13ae: q0 = 16'h00a8; // 0x275c
	13'h13af: q0 = 16'h206d; // 0x275e
	13'h13b0: q0 = 16'h0022; // 0x2760
	13'h13b1: q0 = 16'h3215; // 0x2762
	13'h13b2: q0 = 16'h48c1; // 0x2764
	13'h13b3: q0 = 16'hd2bc; // 0x2766
	13'h13b4: q0 = 16'h0000; // 0x2768
	13'h13b5: q0 = 16'hca18; // 0x276a
	13'h13b6: q0 = 16'h2241; // 0x276c
	13'h13b7: q0 = 16'h1211; // 0x276e
	13'h13b8: q0 = 16'h4881; // 0x2770
	13'h13b9: q0 = 16'hd27c; // 0x2772
	13'h13ba: q0 = 16'h005a; // 0x2774
	13'h13bb: q0 = 16'h3141; // 0x2776
	13'h13bc: q0 = 16'h0004; // 0x2778
	13'h13bd: q0 = 16'h0c55; // 0x277a
	13'h13be: q0 = 16'h0005; // 0x277c
	13'h13bf: q0 = 16'h6f12; // 0x277e
	13'h13c0: q0 = 16'h0c55; // 0x2780
	13'h13c1: q0 = 16'h001f; // 0x2782
	13'h13c2: q0 = 16'h6d06; // 0x2784
	13'h13c3: q0 = 16'h0c55; // 0x2786
	13'h13c4: q0 = 16'h0029; // 0x2788
	13'h13c5: q0 = 16'h6f06; // 0x278a
	13'h13c6: q0 = 16'h0c55; // 0x278c
	13'h13c7: q0 = 16'h0043; // 0x278e
	13'h13c8: q0 = 16'h6d16; // 0x2790
	13'h13c9: q0 = 16'h206d; // 0x2792
	13'h13ca: q0 = 16'h001e; // 0x2794
	13'h13cb: q0 = 16'h317c; // 0x2796
	13'h13cc: q0 = 16'h002c; // 0x2798
	13'h13cd: q0 = 16'h0004; // 0x279a
	13'h13ce: q0 = 16'h302d; // 0x279c
	13'h13cf: q0 = 16'h000e; // 0x279e
	13'h13d0: q0 = 16'h807c; // 0x27a0
	13'h13d1: q0 = 16'h0200; // 0x27a2
	13'h13d2: q0 = 16'h3b40; // 0x27a4
	13'h13d3: q0 = 16'h000e; // 0x27a6
	13'h13d4: q0 = 16'h605a; // 0x27a8
	13'h13d5: q0 = 16'h206d; // 0x27aa
	13'h13d6: q0 = 16'h0022; // 0x27ac
	13'h13d7: q0 = 16'h3215; // 0x27ae
	13'h13d8: q0 = 16'h48c1; // 0x27b0
	13'h13d9: q0 = 16'hd2bc; // 0x27b2
	13'h13da: q0 = 16'h0000; // 0x27b4
	13'h13db: q0 = 16'hca18; // 0x27b6
	13'h13dc: q0 = 16'h2241; // 0x27b8
	13'h13dd: q0 = 16'h1211; // 0x27ba
	13'h13de: q0 = 16'h4881; // 0x27bc
	13'h13df: q0 = 16'hd27c; // 0x27be
	13'h13e0: q0 = 16'h005a; // 0x27c0
	13'h13e1: q0 = 16'h3141; // 0x27c2
	13'h13e2: q0 = 16'h0004; // 0x27c4
	13'h13e3: q0 = 16'h603c; // 0x27c6
	13'h13e4: q0 = 16'h302d; // 0x27c8
	13'h13e5: q0 = 16'h000e; // 0x27ca
	13'h13e6: q0 = 16'h807c; // 0x27cc
	13'h13e7: q0 = 16'h0400; // 0x27ce
	13'h13e8: q0 = 16'h3b40; // 0x27d0
	13'h13e9: q0 = 16'h000e; // 0x27d2
	13'h13ea: q0 = 16'h302d; // 0x27d4
	13'h13eb: q0 = 16'h000e; // 0x27d6
	13'h13ec: q0 = 16'h807c; // 0x27d8
	13'h13ed: q0 = 16'h0100; // 0x27da
	13'h13ee: q0 = 16'h3b40; // 0x27dc
	13'h13ef: q0 = 16'h000e; // 0x27de
	13'h13f0: q0 = 16'h6022; // 0x27e0
	13'h13f1: q0 = 16'h206d; // 0x27e2
	13'h13f2: q0 = 16'h0022; // 0x27e4
	13'h13f3: q0 = 16'h317c; // 0x27e6
	13'h13f4: q0 = 16'h0059; // 0x27e8
	13'h13f5: q0 = 16'h0004; // 0x27ea
	13'h13f6: q0 = 16'h6016; // 0x27ec
	13'h13f7: q0 = 16'h6014; // 0x27ee
	13'h13f8: q0 = 16'hb07c; // 0x27f0
	13'h13f9: q0 = 16'h0007; // 0x27f2
	13'h13fa: q0 = 16'h620e; // 0x27f4
	13'h13fb: q0 = 16'he540; // 0x27f6
	13'h13fc: q0 = 16'h3040; // 0x27f8
	13'h13fd: q0 = 16'hd1fc; // 0x27fa
	13'h13fe: q0 = 16'h0000; // 0x27fc
	13'h13ff: q0 = 16'hc810; // 0x27fe
	13'h1400: q0 = 16'h2050; // 0x2800
	13'h1401: q0 = 16'h4ed0; // 0x2802
	13'h1402: q0 = 16'h082d; // 0x2804
	13'h1403: q0 = 16'h0002; // 0x2806
	13'h1404: q0 = 16'h000e; // 0x2808
	13'h1405: q0 = 16'h6742; // 0x280a
	13'h1406: q0 = 16'h206d; // 0x280c
	13'h1407: q0 = 16'h0026; // 0x280e
	13'h1408: q0 = 16'h226d; // 0x2810
	13'h1409: q0 = 16'h001a; // 0x2812
	13'h140a: q0 = 16'h3211; // 0x2814
	13'h140b: q0 = 16'hd27c; // 0x2816
	13'h140c: q0 = 16'h0031; // 0x2818
	13'h140d: q0 = 16'h5341; // 0x281a
	13'h140e: q0 = 16'h3141; // 0x281c
	13'h140f: q0 = 16'h0004; // 0x281e
	13'h1410: q0 = 16'h3e95; // 0x2820
	13'h1411: q0 = 16'h202d; // 0x2822
	13'h1412: q0 = 16'h0026; // 0x2824
	13'h1413: q0 = 16'h5c80; // 0x2826
	13'h1414: q0 = 16'h2f00; // 0x2828
	13'h1415: q0 = 16'h4eb9; // 0x282a
	13'h1416: q0 = 16'h0000; // 0x282c
	13'h1417: q0 = 16'h3ee6; // 0x282e
	13'h1418: q0 = 16'h4a9f; // 0x2830
	13'h1419: q0 = 16'h206d; // 0x2832
	13'h141a: q0 = 16'h0022; // 0x2834
	13'h141b: q0 = 16'h3215; // 0x2836
	13'h141c: q0 = 16'h48c1; // 0x2838
	13'h141d: q0 = 16'hd2bc; // 0x283a
	13'h141e: q0 = 16'h0000; // 0x283c
	13'h141f: q0 = 16'hca18; // 0x283e
	13'h1420: q0 = 16'h2241; // 0x2840
	13'h1421: q0 = 16'h1211; // 0x2842
	13'h1422: q0 = 16'h4881; // 0x2844
	13'h1423: q0 = 16'hd27c; // 0x2846
	13'h1424: q0 = 16'h005a; // 0x2848
	13'h1425: q0 = 16'h3141; // 0x284a
	13'h1426: q0 = 16'h0004; // 0x284c
	13'h1427: q0 = 16'h082d; // 0x284e
	13'h1428: q0 = 16'h0000; // 0x2850
	13'h1429: q0 = 16'h000e; // 0x2852
	13'h142a: q0 = 16'h6716; // 0x2854
	13'h142b: q0 = 16'h3b7c; // 0x2856
	13'h142c: q0 = 16'h0007; // 0x2858
	13'h142d: q0 = 16'h000c; // 0x285a
	13'h142e: q0 = 16'h206d; // 0x285c
	13'h142f: q0 = 16'h001e; // 0x285e
	13'h1430: q0 = 16'h322d; // 0x2860
	13'h1431: q0 = 16'h0008; // 0x2862
	13'h1432: q0 = 16'hd27c; // 0x2864
	13'h1433: q0 = 16'h0067; // 0x2866
	13'h1434: q0 = 16'h3141; // 0x2868
	13'h1435: q0 = 16'h0004; // 0x286a
	13'h1436: q0 = 16'hbe7c; // 0x286c
	13'h1437: q0 = 16'h0002; // 0x286e
	13'h1438: q0 = 16'h6730; // 0x2870
	13'h1439: q0 = 16'h3039; // 0x2872
	13'h143a: q0 = 16'h0001; // 0x2874
	13'h143b: q0 = 16'h8a76; // 0x2876
	13'h143c: q0 = 16'h226d; // 0x2878
	13'h143d: q0 = 16'h001a; // 0x287a
	13'h143e: q0 = 16'h4281; // 0x287c
	13'h143f: q0 = 16'h3211; // 0x287e
	13'h1440: q0 = 16'he260; // 0x2880
	13'h1441: q0 = 16'hc07c; // 0x2882
	13'h1442: q0 = 16'h0030; // 0x2884
	13'h1443: q0 = 16'h661a; // 0x2886
	13'h1444: q0 = 16'h206d; // 0x2888
	13'h1445: q0 = 16'h0022; // 0x288a
	13'h1446: q0 = 16'h322e; // 0x288c
	13'h1447: q0 = 16'hfff6; // 0x288e
	13'h1448: q0 = 16'h5341; // 0x2890
	13'h1449: q0 = 16'he341; // 0x2892
	13'h144a: q0 = 16'h48c1; // 0x2894
	13'h144b: q0 = 16'hd2bc; // 0x2896
	13'h144c: q0 = 16'h0000; // 0x2898
	13'h144d: q0 = 16'hc802; // 0x289a
	13'h144e: q0 = 16'h2241; // 0x289c
	13'h144f: q0 = 16'h3151; // 0x289e
	13'h1450: q0 = 16'h0006; // 0x28a0
	13'h1451: q0 = 16'h206d; // 0x28a2
	13'h1452: q0 = 16'h001e; // 0x28a4
	13'h1453: q0 = 16'h322e; // 0x28a6
	13'h1454: q0 = 16'hfff6; // 0x28a8
	13'h1455: q0 = 16'h5341; // 0x28aa
	13'h1456: q0 = 16'he341; // 0x28ac
	13'h1457: q0 = 16'h48c1; // 0x28ae
	13'h1458: q0 = 16'hd2bc; // 0x28b0
	13'h1459: q0 = 16'h0000; // 0x28b2
	13'h145a: q0 = 16'hc7f8; // 0x28b4
	13'h145b: q0 = 16'h2241; // 0x28b6
	13'h145c: q0 = 16'h3151; // 0x28b8
	13'h145d: q0 = 16'h0006; // 0x28ba
	13'h145e: q0 = 16'h206d; // 0x28bc
	13'h145f: q0 = 16'h0026; // 0x28be
	13'h1460: q0 = 16'h226d; // 0x28c0
	13'h1461: q0 = 16'h001e; // 0x28c2
	13'h1462: q0 = 16'h3169; // 0x28c4
	13'h1463: q0 = 16'h0006; // 0x28c6
	13'h1464: q0 = 16'h0006; // 0x28c8
	13'h1465: q0 = 16'h3e95; // 0x28ca
	13'h1466: q0 = 16'h202d; // 0x28cc
	13'h1467: q0 = 16'h001e; // 0x28ce
	13'h1468: q0 = 16'h5c80; // 0x28d0
	13'h1469: q0 = 16'h2f00; // 0x28d2
	13'h146a: q0 = 16'h4eb9; // 0x28d4
	13'h146b: q0 = 16'h0000; // 0x28d6
	13'h146c: q0 = 16'h3ee6; // 0x28d8
	13'h146d: q0 = 16'h4a9f; // 0x28da
	13'h146e: q0 = 16'h3e95; // 0x28dc
	13'h146f: q0 = 16'h202d; // 0x28de
	13'h1470: q0 = 16'h0022; // 0x28e0
	13'h1471: q0 = 16'h5c80; // 0x28e2
	13'h1472: q0 = 16'h2f00; // 0x28e4
	13'h1473: q0 = 16'h4eb9; // 0x28e6
	13'h1474: q0 = 16'h0000; // 0x28e8
	13'h1475: q0 = 16'h3ee6; // 0x28ea
	13'h1476: q0 = 16'h4a9f; // 0x28ec
	13'h1477: q0 = 16'h2ebc; // 0x28ee
	13'h1478: q0 = 16'h0000; // 0x28f0
	13'h1479: q0 = 16'hfc54; // 0x28f2
	13'h147a: q0 = 16'h4eb9; // 0x28f4
	13'h147b: q0 = 16'h0000; // 0x28f6
	13'h147c: q0 = 16'h7dd8; // 0x28f8
	13'h147d: q0 = 16'h302d; // 0x28fa
	13'h147e: q0 = 16'h000e; // 0x28fc
	13'h147f: q0 = 16'hc07c; // 0x28fe
	13'h1480: q0 = 16'hfff0; // 0x2900
	13'h1481: q0 = 16'h807c; // 0x2902
	13'h1482: q0 = 16'h0001; // 0x2904
	13'h1483: q0 = 16'h3b40; // 0x2906
	13'h1484: q0 = 16'h000e; // 0x2908
	13'h1485: q0 = 16'h6004; // 0x290a
	13'h1486: q0 = 16'h6002; // 0x290c
	13'h1487: q0 = 16'h60fc; // 0x290e
	13'h1488: q0 = 16'h4a9f; // 0x2910
	13'h1489: q0 = 16'h4cdf; // 0x2912
	13'h148a: q0 = 16'h2080; // 0x2914
	13'h148b: q0 = 16'h4e5e; // 0x2916
	13'h148c: q0 = 16'h4e75; // 0x2918
	13'h148d: q0 = 16'h4e56; // 0x291a
	13'h148e: q0 = 16'h0000; // 0x291c
	13'h148f: q0 = 16'h48e7; // 0x291e
	13'h1490: q0 = 16'h0104; // 0x2920
	13'h1491: q0 = 16'h2a6e; // 0x2922
	13'h1492: q0 = 16'h0008; // 0x2924
	13'h1493: q0 = 16'h302d; // 0x2926
	13'h1494: q0 = 16'h000e; // 0x2928
	13'h1495: q0 = 16'hc07c; // 0x292a
	13'h1496: q0 = 16'h000f; // 0x292c
	13'h1497: q0 = 16'hb07c; // 0x292e
	13'h1498: q0 = 16'h0002; // 0x2930
	13'h1499: q0 = 16'h662c; // 0x2932
	13'h149a: q0 = 16'h4aad; // 0x2934
	13'h149b: q0 = 16'h002a; // 0x2936
	13'h149c: q0 = 16'h6622; // 0x2938
	13'h149d: q0 = 16'h4eb9; // 0x293a
	13'h149e: q0 = 16'h0000; // 0x293c
	13'h149f: q0 = 16'h4ec6; // 0x293e
	13'h14a0: q0 = 16'h4a40; // 0x2940
	13'h14a1: q0 = 16'h6618; // 0x2942
	13'h14a2: q0 = 16'h4eb9; // 0x2944
	13'h14a3: q0 = 16'h0000; // 0x2946
	13'h14a4: q0 = 16'h4738; // 0x2948
	13'h14a5: q0 = 16'hb07c; // 0x294a
	13'h14a6: q0 = 16'h0002; // 0x294c
	13'h14a7: q0 = 16'h670c; // 0x294e
	13'h14a8: q0 = 16'h4257; // 0x2950
	13'h14a9: q0 = 16'h2f0d; // 0x2952
	13'h14aa: q0 = 16'h4eb9; // 0x2954
	13'h14ab: q0 = 16'h0000; // 0x2956
	13'h14ac: q0 = 16'h2c02; // 0x2958
	13'h14ad: q0 = 16'h4a9f; // 0x295a
	13'h14ae: q0 = 16'h6000; // 0x295c
	13'h14af: q0 = 16'h01ae; // 0x295e
	13'h14b0: q0 = 16'h302d; // 0x2960
	13'h14b1: q0 = 16'h000e; // 0x2962
	13'h14b2: q0 = 16'hc07c; // 0x2964
	13'h14b3: q0 = 16'h000f; // 0x2966
	13'h14b4: q0 = 16'hb07c; // 0x2968
	13'h14b5: q0 = 16'h0003; // 0x296a
	13'h14b6: q0 = 16'h6600; // 0x296c
	13'h14b7: q0 = 16'h00a2; // 0x296e
	13'h14b8: q0 = 16'h0c6d; // 0x2970
	13'h14b9: q0 = 16'h000b; // 0x2972
	13'h14ba: q0 = 16'h0008; // 0x2974
	13'h14bb: q0 = 16'h6f0c; // 0x2976
	13'h14bc: q0 = 16'h2e8d; // 0x2978
	13'h14bd: q0 = 16'h4eb9; // 0x297a
	13'h14be: q0 = 16'h0000; // 0x297c
	13'h14bf: q0 = 16'h2ec2; // 0x297e
	13'h14c0: q0 = 16'h6000; // 0x2980
	13'h14c1: q0 = 16'h008a; // 0x2982
	13'h14c2: q0 = 16'h206d; // 0x2984
	13'h14c3: q0 = 16'h001e; // 0x2986
	13'h14c4: q0 = 16'h322d; // 0x2988
	13'h14c5: q0 = 16'h0008; // 0x298a
	13'h14c6: q0 = 16'h5341; // 0x298c
	13'h14c7: q0 = 16'h48c1; // 0x298e
	13'h14c8: q0 = 16'hd2bc; // 0x2990
	13'h14c9: q0 = 16'h0000; // 0x2992
	13'h14ca: q0 = 16'hc884; // 0x2994
	13'h14cb: q0 = 16'h2241; // 0x2996
	13'h14cc: q0 = 16'h1211; // 0x2998
	13'h14cd: q0 = 16'h4881; // 0x299a
	13'h14ce: q0 = 16'h3141; // 0x299c
	13'h14cf: q0 = 16'h0004; // 0x299e
	13'h14d0: q0 = 16'h206d; // 0x29a0
	13'h14d1: q0 = 16'h0022; // 0x29a2
	13'h14d2: q0 = 16'h322d; // 0x29a4
	13'h14d3: q0 = 16'h0008; // 0x29a6
	13'h14d4: q0 = 16'h5341; // 0x29a8
	13'h14d5: q0 = 16'h48c1; // 0x29aa
	13'h14d6: q0 = 16'hd2bc; // 0x29ac
	13'h14d7: q0 = 16'h0000; // 0x29ae
	13'h14d8: q0 = 16'hc890; // 0x29b0
	13'h14d9: q0 = 16'h2241; // 0x29b2
	13'h14da: q0 = 16'h1211; // 0x29b4
	13'h14db: q0 = 16'h4881; // 0x29b6
	13'h14dc: q0 = 16'h3141; // 0x29b8
	13'h14dd: q0 = 16'h0004; // 0x29ba
	13'h14de: q0 = 16'h206d; // 0x29bc
	13'h14df: q0 = 16'h0026; // 0x29be
	13'h14e0: q0 = 16'h226d; // 0x29c0
	13'h14e1: q0 = 16'h001a; // 0x29c2
	13'h14e2: q0 = 16'h3211; // 0x29c4
	13'h14e3: q0 = 16'h5341; // 0x29c6
	13'h14e4: q0 = 16'he541; // 0x29c8
	13'h14e5: q0 = 16'h48c1; // 0x29ca
	13'h14e6: q0 = 16'hd2bc; // 0x29cc
	13'h14e7: q0 = 16'h0001; // 0x29ce
	13'h14e8: q0 = 16'h85fe; // 0x29d0
	13'h14e9: q0 = 16'h2241; // 0x29d2
	13'h14ea: q0 = 16'h2211; // 0x29d4
	13'h14eb: q0 = 16'h342d; // 0x29d6
	13'h14ec: q0 = 16'h0008; // 0x29d8
	13'h14ed: q0 = 16'h5342; // 0x29da
	13'h14ee: q0 = 16'h48c2; // 0x29dc
	13'h14ef: q0 = 16'hd282; // 0x29de
	13'h14f0: q0 = 16'h2241; // 0x29e0
	13'h14f1: q0 = 16'h1211; // 0x29e2
	13'h14f2: q0 = 16'h4881; // 0x29e4
	13'h14f3: q0 = 16'h3141; // 0x29e6
	13'h14f4: q0 = 16'h0004; // 0x29e8
	13'h14f5: q0 = 16'h3ead; // 0x29ea
	13'h14f6: q0 = 16'h0018; // 0x29ec
	13'h14f7: q0 = 16'h302d; // 0x29ee
	13'h14f8: q0 = 16'h0008; // 0x29f0
	13'h14f9: q0 = 16'h5340; // 0x29f2
	13'h14fa: q0 = 16'he140; // 0x29f4
	13'h14fb: q0 = 16'h9157; // 0x29f6
	13'h14fc: q0 = 16'h206d; // 0x29f8
	13'h14fd: q0 = 16'h001e; // 0x29fa
	13'h14fe: q0 = 16'h3f10; // 0x29fc
	13'h14ff: q0 = 16'h2f0d; // 0x29fe
	13'h1500: q0 = 16'h4eb9; // 0x2a00
	13'h1501: q0 = 16'h0000; // 0x2a02
	13'h1502: q0 = 16'h2dc2; // 0x2a04
	13'h1503: q0 = 16'h5c4f; // 0x2a06
	13'h1504: q0 = 16'h526d; // 0x2a08
	13'h1505: q0 = 16'h0008; // 0x2a0a
	13'h1506: q0 = 16'h6000; // 0x2a0c
	13'h1507: q0 = 16'h00fe; // 0x2a0e
	13'h1508: q0 = 16'h302d; // 0x2a10
	13'h1509: q0 = 16'h000e; // 0x2a12
	13'h150a: q0 = 16'hc07c; // 0x2a14
	13'h150b: q0 = 16'h000f; // 0x2a16
	13'h150c: q0 = 16'hb07c; // 0x2a18
	13'h150d: q0 = 16'h0004; // 0x2a1a
	13'h150e: q0 = 16'h6600; // 0x2a1c
	13'h150f: q0 = 16'h00ea; // 0x2a1e
	13'h1510: q0 = 16'h0c6d; // 0x2a20
	13'h1511: q0 = 16'h000b; // 0x2a22
	13'h1512: q0 = 16'h0008; // 0x2a24
	13'h1513: q0 = 16'h6f14; // 0x2a26
	13'h1514: q0 = 16'h4a79; // 0x2a28
	13'h1515: q0 = 16'h0001; // 0x2a2a
	13'h1516: q0 = 16'h7b9e; // 0x2a2c
	13'h1517: q0 = 16'h6608; // 0x2a2e
	13'h1518: q0 = 16'h2e8d; // 0x2a30
	13'h1519: q0 = 16'h4eb9; // 0x2a32
	13'h151a: q0 = 16'h0000; // 0x2a34
	13'h151b: q0 = 16'h1f50; // 0x2a36
	13'h151c: q0 = 16'h6000; // 0x2a38
	13'h151d: q0 = 16'h00d2; // 0x2a3a
	13'h151e: q0 = 16'h206d; // 0x2a3c
	13'h151f: q0 = 16'h001e; // 0x2a3e
	13'h1520: q0 = 16'h720b; // 0x2a40
	13'h1521: q0 = 16'h926d; // 0x2a42
	13'h1522: q0 = 16'h0008; // 0x2a44
	13'h1523: q0 = 16'h48c1; // 0x2a46
	13'h1524: q0 = 16'hd2bc; // 0x2a48
	13'h1525: q0 = 16'h0000; // 0x2a4a
	13'h1526: q0 = 16'hc884; // 0x2a4c
	13'h1527: q0 = 16'h2241; // 0x2a4e
	13'h1528: q0 = 16'h1211; // 0x2a50
	13'h1529: q0 = 16'h4881; // 0x2a52
	13'h152a: q0 = 16'h3141; // 0x2a54
	13'h152b: q0 = 16'h0004; // 0x2a56
	13'h152c: q0 = 16'h206d; // 0x2a58
	13'h152d: q0 = 16'h0022; // 0x2a5a
	13'h152e: q0 = 16'h720b; // 0x2a5c
	13'h152f: q0 = 16'h926d; // 0x2a5e
	13'h1530: q0 = 16'h0008; // 0x2a60
	13'h1531: q0 = 16'h48c1; // 0x2a62
	13'h1532: q0 = 16'hd2bc; // 0x2a64
	13'h1533: q0 = 16'h0000; // 0x2a66
	13'h1534: q0 = 16'hc890; // 0x2a68
	13'h1535: q0 = 16'h2241; // 0x2a6a
	13'h1536: q0 = 16'h1211; // 0x2a6c
	13'h1537: q0 = 16'h4881; // 0x2a6e
	13'h1538: q0 = 16'h3141; // 0x2a70
	13'h1539: q0 = 16'h0004; // 0x2a72
	13'h153a: q0 = 16'h206d; // 0x2a74
	13'h153b: q0 = 16'h0026; // 0x2a76
	13'h153c: q0 = 16'h226d; // 0x2a78
	13'h153d: q0 = 16'h001a; // 0x2a7a
	13'h153e: q0 = 16'h3211; // 0x2a7c
	13'h153f: q0 = 16'h5341; // 0x2a7e
	13'h1540: q0 = 16'he541; // 0x2a80
	13'h1541: q0 = 16'h48c1; // 0x2a82
	13'h1542: q0 = 16'hd2bc; // 0x2a84
	13'h1543: q0 = 16'h0001; // 0x2a86
	13'h1544: q0 = 16'h85fe; // 0x2a88
	13'h1545: q0 = 16'h2241; // 0x2a8a
	13'h1546: q0 = 16'h2211; // 0x2a8c
	13'h1547: q0 = 16'hd2bc; // 0x2a8e
	13'h1548: q0 = 16'h0000; // 0x2a90
	13'h1549: q0 = 16'h000b; // 0x2a92
	13'h154a: q0 = 16'h342d; // 0x2a94
	13'h154b: q0 = 16'h0008; // 0x2a96
	13'h154c: q0 = 16'h48c2; // 0x2a98
	13'h154d: q0 = 16'h9282; // 0x2a9a
	13'h154e: q0 = 16'h2241; // 0x2a9c
	13'h154f: q0 = 16'h1211; // 0x2a9e
	13'h1550: q0 = 16'h4881; // 0x2aa0
	13'h1551: q0 = 16'h3141; // 0x2aa2
	13'h1552: q0 = 16'h0004; // 0x2aa4
	13'h1553: q0 = 16'h3ead; // 0x2aa6
	13'h1554: q0 = 16'h0018; // 0x2aa8
	13'h1555: q0 = 16'h700b; // 0x2aaa
	13'h1556: q0 = 16'h906d; // 0x2aac
	13'h1557: q0 = 16'h0008; // 0x2aae
	13'h1558: q0 = 16'he140; // 0x2ab0
	13'h1559: q0 = 16'h9157; // 0x2ab2
	13'h155a: q0 = 16'h206d; // 0x2ab4
	13'h155b: q0 = 16'h001e; // 0x2ab6
	13'h155c: q0 = 16'h3f10; // 0x2ab8
	13'h155d: q0 = 16'h2f0d; // 0x2aba
	13'h155e: q0 = 16'h4eb9; // 0x2abc
	13'h155f: q0 = 16'h0000; // 0x2abe
	13'h1560: q0 = 16'h2dc2; // 0x2ac0
	13'h1561: q0 = 16'h5c4f; // 0x2ac2
	13'h1562: q0 = 16'h4a6d; // 0x2ac4
	13'h1563: q0 = 16'h000a; // 0x2ac6
	13'h1564: q0 = 16'h6638; // 0x2ac8
	13'h1565: q0 = 16'h3b6d; // 0x2aca
	13'h1566: q0 = 16'h000c; // 0x2acc
	13'h1567: q0 = 16'h000a; // 0x2ace
	13'h1568: q0 = 16'h526d; // 0x2ad0
	13'h1569: q0 = 16'h0008; // 0x2ad2
	13'h156a: q0 = 16'h0c6d; // 0x2ad4
	13'h156b: q0 = 16'h0002; // 0x2ad6
	13'h156c: q0 = 16'h0008; // 0x2ad8
	13'h156d: q0 = 16'h6624; // 0x2ada
	13'h156e: q0 = 16'h4a79; // 0x2adc
	13'h156f: q0 = 16'h0001; // 0x2ade
	13'h1570: q0 = 16'h8676; // 0x2ae0
	13'h1571: q0 = 16'h661c; // 0x2ae2
	13'h1572: q0 = 16'h206d; // 0x2ae4
	13'h1573: q0 = 16'h001a; // 0x2ae6
	13'h1574: q0 = 16'h3010; // 0x2ae8
	13'h1575: q0 = 16'h5340; // 0x2aea
	13'h1576: q0 = 16'he540; // 0x2aec
	13'h1577: q0 = 16'h48c0; // 0x2aee
	13'h1578: q0 = 16'hd0bc; // 0x2af0
	13'h1579: q0 = 16'h0000; // 0x2af2
	13'h157a: q0 = 16'hc830; // 0x2af4
	13'h157b: q0 = 16'h2040; // 0x2af6
	13'h157c: q0 = 16'h2e90; // 0x2af8
	13'h157d: q0 = 16'h4eb9; // 0x2afa
	13'h157e: q0 = 16'h0000; // 0x2afc
	13'h157f: q0 = 16'h7dd8; // 0x2afe
	13'h1580: q0 = 16'h6004; // 0x2b00
	13'h1581: q0 = 16'h536d; // 0x2b02
	13'h1582: q0 = 16'h000a; // 0x2b04
	13'h1583: q0 = 16'h6004; // 0x2b06
	13'h1584: q0 = 16'h6002; // 0x2b08
	13'h1585: q0 = 16'h60fc; // 0x2b0a
	13'h1586: q0 = 16'h4a9f; // 0x2b0c
	13'h1587: q0 = 16'h4cdf; // 0x2b0e
	13'h1588: q0 = 16'h2000; // 0x2b10
	13'h1589: q0 = 16'h4e5e; // 0x2b12
	13'h158a: q0 = 16'h4e75; // 0x2b14
	13'h158b: q0 = 16'h4e56; // 0x2b16
	13'h158c: q0 = 16'hfffc; // 0x2b18
	13'h158d: q0 = 16'h48e7; // 0x2b1a
	13'h158e: q0 = 16'h3f00; // 0x2b1c
	13'h158f: q0 = 16'h4eb9; // 0x2b1e
	13'h1590: q0 = 16'h0000; // 0x2b20
	13'h1591: q0 = 16'h4ee2; // 0x2b22
	13'h1592: q0 = 16'h3800; // 0x2b24
	13'h1593: q0 = 16'h4eb9; // 0x2b26
	13'h1594: q0 = 16'h0000; // 0x2b28
	13'h1595: q0 = 16'h4f30; // 0x2b2a
	13'h1596: q0 = 16'h3600; // 0x2b2c
	13'h1597: q0 = 16'h4eb9; // 0x2b2e
	13'h1598: q0 = 16'h0000; // 0x2b30
	13'h1599: q0 = 16'h4f00; // 0x2b32
	13'h159a: q0 = 16'h3d40; // 0x2b34
	13'h159b: q0 = 16'hfffe; // 0x2b36
	13'h159c: q0 = 16'h4eb9; // 0x2b38
	13'h159d: q0 = 16'h0000; // 0x2b3a
	13'h159e: q0 = 16'h4f50; // 0x2b3c
	13'h159f: q0 = 16'h3d40; // 0x2b3e
	13'h15a0: q0 = 16'hfffc; // 0x2b40
	13'h15a1: q0 = 16'h3a2e; // 0x2b42
	13'h15a2: q0 = 16'h0008; // 0x2b44
	13'h15a3: q0 = 16'h4a6e; // 0x2b46
	13'h15a4: q0 = 16'hfffe; // 0x2b48
	13'h15a5: q0 = 16'h6608; // 0x2b4a
	13'h15a6: q0 = 16'h4a6e; // 0x2b4c
	13'h15a7: q0 = 16'hfffc; // 0x2b4e
	13'h15a8: q0 = 16'h6602; // 0x2b50
	13'h15a9: q0 = 16'h7a01; // 0x2b52
	13'h15aa: q0 = 16'h3005; // 0x2b54
	13'h15ab: q0 = 16'h6056; // 0x2b56
	13'h15ac: q0 = 16'h3c03; // 0x2b58
	13'h15ad: q0 = 16'h3e04; // 0x2b5a
	13'h15ae: q0 = 16'h6066; // 0x2b5c
	13'h15af: q0 = 16'h3c03; // 0x2b5e
	13'h15b0: q0 = 16'h9c79; // 0x2b60
	13'h15b1: q0 = 16'h0001; // 0x2b62
	13'h15b2: q0 = 16'h8938; // 0x2b64
	13'h15b3: q0 = 16'he246; // 0x2b66
	13'h15b4: q0 = 16'hdc79; // 0x2b68
	13'h15b5: q0 = 16'h0001; // 0x2b6a
	13'h15b6: q0 = 16'h8938; // 0x2b6c
	13'h15b7: q0 = 16'h3e04; // 0x2b6e
	13'h15b8: q0 = 16'h9e79; // 0x2b70
	13'h15b9: q0 = 16'h0001; // 0x2b72
	13'h15ba: q0 = 16'h8936; // 0x2b74
	13'h15bb: q0 = 16'he247; // 0x2b76
	13'h15bc: q0 = 16'hde79; // 0x2b78
	13'h15bd: q0 = 16'h0001; // 0x2b7a
	13'h15be: q0 = 16'h8936; // 0x2b7c
	13'h15bf: q0 = 16'h6044; // 0x2b7e
	13'h15c0: q0 = 16'h3c2e; // 0x2b80
	13'h15c1: q0 = 16'hfffc; // 0x2b82
	13'h15c2: q0 = 16'he946; // 0x2b84
	13'h15c3: q0 = 16'hdc43; // 0x2b86
	13'h15c4: q0 = 16'h3e2e; // 0x2b88
	13'h15c5: q0 = 16'hfffe; // 0x2b8a
	13'h15c6: q0 = 16'he947; // 0x2b8c
	13'h15c7: q0 = 16'hde44; // 0x2b8e
	13'h15c8: q0 = 16'h6032; // 0x2b90
	13'h15c9: q0 = 16'h3003; // 0x2b92
	13'h15ca: q0 = 16'h322e; // 0x2b94
	13'h15cb: q0 = 16'hfffc; // 0x2b96
	13'h15cc: q0 = 16'he941; // 0x2b98
	13'h15cd: q0 = 16'h9041; // 0x2b9a
	13'h15ce: q0 = 16'h3c00; // 0x2b9c
	13'h15cf: q0 = 16'h3004; // 0x2b9e
	13'h15d0: q0 = 16'h322e; // 0x2ba0
	13'h15d1: q0 = 16'hfffe; // 0x2ba2
	13'h15d2: q0 = 16'he941; // 0x2ba4
	13'h15d3: q0 = 16'h9041; // 0x2ba6
	13'h15d4: q0 = 16'h3e00; // 0x2ba8
	13'h15d5: q0 = 16'h6018; // 0x2baa
	13'h15d6: q0 = 16'h6016; // 0x2bac
	13'h15d7: q0 = 16'h5340; // 0x2bae
	13'h15d8: q0 = 16'hb07c; // 0x2bb0
	13'h15d9: q0 = 16'h0003; // 0x2bb2
	13'h15da: q0 = 16'h620e; // 0x2bb4
	13'h15db: q0 = 16'he540; // 0x2bb6
	13'h15dc: q0 = 16'h3040; // 0x2bb8
	13'h15dd: q0 = 16'hd1fc; // 0x2bba
	13'h15de: q0 = 16'h0000; // 0x2bbc
	13'h15df: q0 = 16'hc840; // 0x2bbe
	13'h15e0: q0 = 16'h2050; // 0x2bc0
	13'h15e1: q0 = 16'h4ed0; // 0x2bc2
	13'h15e2: q0 = 16'hbc7c; // 0x2bc4
	13'h15e3: q0 = 16'h1400; // 0x2bc6
	13'h15e4: q0 = 16'h6d06; // 0x2bc8
	13'h15e5: q0 = 16'hbc7c; // 0x2bca
	13'h15e6: q0 = 16'h7400; // 0x2bcc
	13'h15e7: q0 = 16'h6f02; // 0x2bce
	13'h15e8: q0 = 16'h3c03; // 0x2bd0
	13'h15e9: q0 = 16'hbe7c; // 0x2bd2
	13'h15ea: q0 = 16'h0180; // 0x2bd4
	13'h15eb: q0 = 16'h6d06; // 0x2bd6
	13'h15ec: q0 = 16'hbe7c; // 0x2bd8
	13'h15ed: q0 = 16'h7780; // 0x2bda
	13'h15ee: q0 = 16'h6f02; // 0x2bdc
	13'h15ef: q0 = 16'h3e04; // 0x2bde
	13'h15f0: q0 = 16'h3e86; // 0x2be0
	13'h15f1: q0 = 16'h302e; // 0x2be2
	13'h15f2: q0 = 16'h000c; // 0x2be4
	13'h15f3: q0 = 16'h9157; // 0x2be6
	13'h15f4: q0 = 16'h3f07; // 0x2be8
	13'h15f5: q0 = 16'h302e; // 0x2bea
	13'h15f6: q0 = 16'h000a; // 0x2bec
	13'h15f7: q0 = 16'h9157; // 0x2bee
	13'h15f8: q0 = 16'h4eb9; // 0x2bf0
	13'h15f9: q0 = 16'h0000; // 0x2bf2
	13'h15fa: q0 = 16'h0a1c; // 0x2bf4
	13'h15fb: q0 = 16'h4a5f; // 0x2bf6
	13'h15fc: q0 = 16'h4a9f; // 0x2bf8
	13'h15fd: q0 = 16'h4cdf; // 0x2bfa
	13'h15fe: q0 = 16'h00f8; // 0x2bfc
	13'h15ff: q0 = 16'h4e5e; // 0x2bfe
	13'h1600: q0 = 16'h4e75; // 0x2c00
	13'h1601: q0 = 16'h4e56; // 0x2c02
	13'h1602: q0 = 16'hfffc; // 0x2c04
	13'h1603: q0 = 16'h48e7; // 0x2c06
	13'h1604: q0 = 16'h0104; // 0x2c08
	13'h1605: q0 = 16'h2a6e; // 0x2c0a
	13'h1606: q0 = 16'h0008; // 0x2c0c
	13'h1607: q0 = 16'h3eae; // 0x2c0e
	13'h1608: q0 = 16'h000c; // 0x2c10
	13'h1609: q0 = 16'h200e; // 0x2c12
	13'h160a: q0 = 16'hd0bc; // 0x2c14
	13'h160b: q0 = 16'hffff; // 0x2c16
	13'h160c: q0 = 16'hfffc; // 0x2c18
	13'h160d: q0 = 16'h2f00; // 0x2c1a
	13'h160e: q0 = 16'h200e; // 0x2c1c
	13'h160f: q0 = 16'hd0bc; // 0x2c1e
	13'h1610: q0 = 16'hffff; // 0x2c20
	13'h1611: q0 = 16'hfffe; // 0x2c22
	13'h1612: q0 = 16'h2f00; // 0x2c24
	13'h1613: q0 = 16'h4eb9; // 0x2c26
	13'h1614: q0 = 16'h0000; // 0x2c28
	13'h1615: q0 = 16'h5e3a; // 0x2c2a
	13'h1616: q0 = 16'hbf8f; // 0x2c2c
	13'h1617: q0 = 16'h3eae; // 0x2c2e
	13'h1618: q0 = 16'hfffc; // 0x2c30
	13'h1619: q0 = 16'h3f2e; // 0x2c32
	13'h161a: q0 = 16'hfffe; // 0x2c34
	13'h161b: q0 = 16'h2f0d; // 0x2c36
	13'h161c: q0 = 16'h4eb9; // 0x2c38
	13'h161d: q0 = 16'h0000; // 0x2c3a
	13'h161e: q0 = 16'h2dc2; // 0x2c3c
	13'h161f: q0 = 16'h5c4f; // 0x2c3e
	13'h1620: q0 = 16'h3b6e; // 0x2c40
	13'h1621: q0 = 16'hfffc; // 0x2c42
	13'h1622: q0 = 16'h0018; // 0x2c44
	13'h1623: q0 = 16'h206d; // 0x2c46
	13'h1624: q0 = 16'h001e; // 0x2c48
	13'h1625: q0 = 16'h317c; // 0x2c4a
	13'h1626: q0 = 16'h0017; // 0x2c4c
	13'h1627: q0 = 16'h0006; // 0x2c4e
	13'h1628: q0 = 16'h206d; // 0x2c50
	13'h1629: q0 = 16'h0022; // 0x2c52
	13'h162a: q0 = 16'h317c; // 0x2c54
	13'h162b: q0 = 16'h0008; // 0x2c56
	13'h162c: q0 = 16'h0006; // 0x2c58
	13'h162d: q0 = 16'h206d; // 0x2c5a
	13'h162e: q0 = 16'h0026; // 0x2c5c
	13'h162f: q0 = 16'h317c; // 0x2c5e
	13'h1630: q0 = 16'h0017; // 0x2c60
	13'h1631: q0 = 16'h0006; // 0x2c62
	13'h1632: q0 = 16'h3e95; // 0x2c64
	13'h1633: q0 = 16'h202d; // 0x2c66
	13'h1634: q0 = 16'h001e; // 0x2c68
	13'h1635: q0 = 16'h5c80; // 0x2c6a
	13'h1636: q0 = 16'h2f00; // 0x2c6c
	13'h1637: q0 = 16'h4eb9; // 0x2c6e
	13'h1638: q0 = 16'h0000; // 0x2c70
	13'h1639: q0 = 16'h3ee6; // 0x2c72
	13'h163a: q0 = 16'h4a9f; // 0x2c74
	13'h163b: q0 = 16'h3e95; // 0x2c76
	13'h163c: q0 = 16'h202d; // 0x2c78
	13'h163d: q0 = 16'h0022; // 0x2c7a
	13'h163e: q0 = 16'h5c80; // 0x2c7c
	13'h163f: q0 = 16'h2f00; // 0x2c7e
	13'h1640: q0 = 16'h4eb9; // 0x2c80
	13'h1641: q0 = 16'h0000; // 0x2c82
	13'h1642: q0 = 16'h3ee6; // 0x2c84
	13'h1643: q0 = 16'h4a9f; // 0x2c86
	13'h1644: q0 = 16'h3b7c; // 0x2c88
	13'h1645: q0 = 16'h0001; // 0x2c8a
	13'h1646: q0 = 16'h0008; // 0x2c8c
	13'h1647: q0 = 16'h3b7c; // 0x2c8e
	13'h1648: q0 = 16'h0001; // 0x2c90
	13'h1649: q0 = 16'h000c; // 0x2c92
	13'h164a: q0 = 16'h3b6d; // 0x2c94
	13'h164b: q0 = 16'h000c; // 0x2c96
	13'h164c: q0 = 16'h000a; // 0x2c98
	13'h164d: q0 = 16'h302d; // 0x2c9a
	13'h164e: q0 = 16'h000e; // 0x2c9c
	13'h164f: q0 = 16'hc07c; // 0x2c9e
	13'h1650: q0 = 16'hf0f0; // 0x2ca0
	13'h1651: q0 = 16'h807c; // 0x2ca2
	13'h1652: q0 = 16'h0004; // 0x2ca4
	13'h1653: q0 = 16'h3b40; // 0x2ca6
	13'h1654: q0 = 16'h000e; // 0x2ca8
	13'h1655: q0 = 16'h5279; // 0x2caa
	13'h1656: q0 = 16'h0001; // 0x2cac
	13'h1657: q0 = 16'h86d4; // 0x2cae
	13'h1658: q0 = 16'h4a9f; // 0x2cb0
	13'h1659: q0 = 16'h4cdf; // 0x2cb2
	13'h165a: q0 = 16'h2000; // 0x2cb4
	13'h165b: q0 = 16'h4e5e; // 0x2cb6
	13'h165c: q0 = 16'h4e75; // 0x2cb8
	13'h165d: q0 = 16'h4e56; // 0x2cba
	13'h165e: q0 = 16'h0000; // 0x2cbc
	13'h165f: q0 = 16'h48e7; // 0x2cbe
	13'h1660: q0 = 16'h1f04; // 0x2cc0
	13'h1661: q0 = 16'h4eb9; // 0x2cc2
	13'h1662: q0 = 16'h0000; // 0x2cc4
	13'h1663: q0 = 16'h1e8a; // 0x2cc6
	13'h1664: q0 = 16'h2079; // 0x2cc8
	13'h1665: q0 = 16'h0001; // 0x2cca
	13'h1666: q0 = 16'h7fb8; // 0x2ccc
	13'h1667: q0 = 16'h3010; // 0x2cce
	13'h1668: q0 = 16'h5240; // 0x2cd0
	13'h1669: q0 = 16'h33c0; // 0x2cd2
	13'h166a: q0 = 16'h0001; // 0x2cd4
	13'h166b: q0 = 16'h7fbc; // 0x2cd6
	13'h166c: q0 = 16'h0c79; // 0x2cd8
	13'h166d: q0 = 16'h0004; // 0x2cda
	13'h166e: q0 = 16'h0001; // 0x2cdc
	13'h166f: q0 = 16'h7fbc; // 0x2cde
	13'h1670: q0 = 16'h6f08; // 0x2ce0
	13'h1671: q0 = 16'h33fc; // 0x2ce2
	13'h1672: q0 = 16'h0004; // 0x2ce4
	13'h1673: q0 = 16'h0001; // 0x2ce6
	13'h1674: q0 = 16'h7fbc; // 0x2ce8
	13'h1675: q0 = 16'h3039; // 0x2cea
	13'h1676: q0 = 16'h0001; // 0x2cec
	13'h1677: q0 = 16'h757e; // 0x2cee
	13'h1678: q0 = 16'h5340; // 0x2cf0
	13'h1679: q0 = 16'he340; // 0x2cf2
	13'h167a: q0 = 16'h48c0; // 0x2cf4
	13'h167b: q0 = 16'hd0bc; // 0x2cf6
	13'h167c: q0 = 16'h0000; // 0x2cf8
	13'h167d: q0 = 16'hc8c8; // 0x2cfa
	13'h167e: q0 = 16'h2040; // 0x2cfc
	13'h167f: q0 = 16'h3a10; // 0x2cfe
	13'h1680: q0 = 16'h2079; // 0x2d00
	13'h1681: q0 = 16'h0001; // 0x2d02
	13'h1682: q0 = 16'h7fb8; // 0x2d04
	13'h1683: q0 = 16'h3c10; // 0x2d06
	13'h1684: q0 = 16'hbc7c; // 0x2d08
	13'h1685: q0 = 16'h0003; // 0x2d0a
	13'h1686: q0 = 16'h6e10; // 0x2d0c
	13'h1687: q0 = 16'h7041; // 0x2d0e
	13'h1688: q0 = 16'h3206; // 0x2d10
	13'h1689: q0 = 16'he541; // 0x2d12
	13'h168a: q0 = 16'h9041; // 0x2d14
	13'h168b: q0 = 16'h33c0; // 0x2d16
	13'h168c: q0 = 16'h0001; // 0x2d18
	13'h168d: q0 = 16'h7f28; // 0x2d1a
	13'h168e: q0 = 16'h6030; // 0x2d1c
	13'h168f: q0 = 16'hbc45; // 0x2d1e
	13'h1690: q0 = 16'h6d08; // 0x2d20
	13'h1691: q0 = 16'h4279; // 0x2d22
	13'h1692: q0 = 16'h0001; // 0x2d24
	13'h1693: q0 = 16'h7f28; // 0x2d26
	13'h1694: q0 = 16'h6024; // 0x2d28
	13'h1695: q0 = 16'h7835; // 0x2d2a
	13'h1696: q0 = 16'h3005; // 0x2d2c
	13'h1697: q0 = 16'h5740; // 0x2d2e
	13'h1698: q0 = 16'he240; // 0x2d30
	13'h1699: q0 = 16'hd044; // 0x2d32
	13'h169a: q0 = 16'h48c0; // 0x2d34
	13'h169b: q0 = 16'h3205; // 0x2d36
	13'h169c: q0 = 16'h5741; // 0x2d38
	13'h169d: q0 = 16'h81c1; // 0x2d3a
	13'h169e: q0 = 16'h3206; // 0x2d3c
	13'h169f: q0 = 16'h5741; // 0x2d3e
	13'h16a0: q0 = 16'hc1c1; // 0x2d40
	13'h16a1: q0 = 16'h3f00; // 0x2d42
	13'h16a2: q0 = 16'h3004; // 0x2d44
	13'h16a3: q0 = 16'h905f; // 0x2d46
	13'h16a4: q0 = 16'h33c0; // 0x2d48
	13'h16a5: q0 = 16'h0001; // 0x2d4a
	13'h16a6: q0 = 16'h7f28; // 0x2d4c
	13'h16a7: q0 = 16'h2a7c; // 0x2d4e
	13'h16a8: q0 = 16'h0001; // 0x2d50
	13'h16a9: q0 = 16'h89be; // 0x2d52
	13'h16aa: q0 = 16'h4247; // 0x2d54
	13'h16ab: q0 = 16'hbe79; // 0x2d56
	13'h16ac: q0 = 16'h0001; // 0x2d58
	13'h16ad: q0 = 16'h7fbc; // 0x2d5a
	13'h16ae: q0 = 16'h6c5a; // 0x2d5c
	13'h16af: q0 = 16'h426d; // 0x2d5e
	13'h16b0: q0 = 16'h000e; // 0x2d60
	13'h16b1: q0 = 16'h4255; // 0x2d62
	13'h16b2: q0 = 16'h42ad; // 0x2d64
	13'h16b3: q0 = 16'h0010; // 0x2d66
	13'h16b4: q0 = 16'h3007; // 0x2d68
	13'h16b5: q0 = 16'hc1fc; // 0x2d6a
	13'h16b6: q0 = 16'h0006; // 0x2d6c
	13'h16b7: q0 = 16'hd0bc; // 0x2d6e
	13'h16b8: q0 = 16'h0000; // 0x2d70
	13'h16b9: q0 = 16'hc850; // 0x2d72
	13'h16ba: q0 = 16'h2b40; // 0x2d74
	13'h16bb: q0 = 16'h001a; // 0x2d76
	13'h16bc: q0 = 16'h206d; // 0x2d78
	13'h16bd: q0 = 16'h001a; // 0x2d7a
	13'h16be: q0 = 16'h3010; // 0x2d7c
	13'h16bf: q0 = 16'h5340; // 0x2d7e
	13'h16c0: q0 = 16'hc1fc; // 0x2d80
	13'h16c1: q0 = 16'h000b; // 0x2d82
	13'h16c2: q0 = 16'h48c0; // 0x2d84
	13'h16c3: q0 = 16'hd0bc; // 0x2d86
	13'h16c4: q0 = 16'h0000; // 0x2d88
	13'h16c5: q0 = 16'hc89c; // 0x2d8a
	13'h16c6: q0 = 16'h226d; // 0x2d8c
	13'h16c7: q0 = 16'h001a; // 0x2d8e
	13'h16c8: q0 = 16'h3211; // 0x2d90
	13'h16c9: q0 = 16'h5341; // 0x2d92
	13'h16ca: q0 = 16'he541; // 0x2d94
	13'h16cb: q0 = 16'h48c1; // 0x2d96
	13'h16cc: q0 = 16'hd2bc; // 0x2d98
	13'h16cd: q0 = 16'h0001; // 0x2d9a
	13'h16ce: q0 = 16'h85fe; // 0x2d9c
	13'h16cf: q0 = 16'h2241; // 0x2d9e
	13'h16d0: q0 = 16'h2280; // 0x2da0
	13'h16d1: q0 = 16'h4257; // 0x2da2
	13'h16d2: q0 = 16'h2f0d; // 0x2da4
	13'h16d3: q0 = 16'h4eb9; // 0x2da6
	13'h16d4: q0 = 16'h0000; // 0x2da8
	13'h16d5: q0 = 16'h2c02; // 0x2daa
	13'h16d6: q0 = 16'h4a9f; // 0x2dac
	13'h16d7: q0 = 16'hdbfc; // 0x2dae
	13'h16d8: q0 = 16'h0000; // 0x2db0
	13'h16d9: q0 = 16'h002e; // 0x2db2
	13'h16da: q0 = 16'h5247; // 0x2db4
	13'h16db: q0 = 16'h609e; // 0x2db6
	13'h16dc: q0 = 16'h4a9f; // 0x2db8
	13'h16dd: q0 = 16'h4cdf; // 0x2dba
	13'h16de: q0 = 16'h20f0; // 0x2dbc
	13'h16df: q0 = 16'h4e5e; // 0x2dbe
	13'h16e0: q0 = 16'h4e75; // 0x2dc0
	13'h16e1: q0 = 16'h4e56; // 0x2dc2
	13'h16e2: q0 = 16'h0000; // 0x2dc4
	13'h16e3: q0 = 16'h48e7; // 0x2dc6
	13'h16e4: q0 = 16'h0704; // 0x2dc8
	13'h16e5: q0 = 16'h2a6e; // 0x2dca
	13'h16e6: q0 = 16'h0008; // 0x2dcc
	13'h16e7: q0 = 16'h3e2e; // 0x2dce
	13'h16e8: q0 = 16'h000c; // 0x2dd0
	13'h16e9: q0 = 16'h3c2e; // 0x2dd2
	13'h16ea: q0 = 16'h000e; // 0x2dd4
	13'h16eb: q0 = 16'h206d; // 0x2dd6
	13'h16ec: q0 = 16'h001e; // 0x2dd8
	13'h16ed: q0 = 16'h3087; // 0x2dda
	13'h16ee: q0 = 16'h206d; // 0x2ddc
	13'h16ef: q0 = 16'h001e; // 0x2dde
	13'h16f0: q0 = 16'h3146; // 0x2de0
	13'h16f1: q0 = 16'h0002; // 0x2de2
	13'h16f2: q0 = 16'h206d; // 0x2de4
	13'h16f3: q0 = 16'h0022; // 0x2de6
	13'h16f4: q0 = 16'h3087; // 0x2de8
	13'h16f5: q0 = 16'h082d; // 0x2dea
	13'h16f6: q0 = 16'h0000; // 0x2dec
	13'h16f7: q0 = 16'h000e; // 0x2dee
	13'h16f8: q0 = 16'h6742; // 0x2df0
	13'h16f9: q0 = 16'h0c6d; // 0x2df2
	13'h16fa: q0 = 16'h0012; // 0x2df4
	13'h16fb: q0 = 16'h0008; // 0x2df6
	13'h16fc: q0 = 16'h6f22; // 0x2df8
	13'h16fd: q0 = 16'h0c6d; // 0x2dfa
	13'h16fe: q0 = 16'h0036; // 0x2dfc
	13'h16ff: q0 = 16'h0008; // 0x2dfe
	13'h1700: q0 = 16'h6e1a; // 0x2e00
	13'h1701: q0 = 16'h0c55; // 0x2e02
	13'h1702: q0 = 16'h0012; // 0x2e04
	13'h1703: q0 = 16'h6f06; // 0x2e06
	13'h1704: q0 = 16'h0c55; // 0x2e08
	13'h1705: q0 = 16'h0036; // 0x2e0a
	13'h1706: q0 = 16'h6f0c; // 0x2e0c
	13'h1707: q0 = 16'h206d; // 0x2e0e
	13'h1708: q0 = 16'h0022; // 0x2e10
	13'h1709: q0 = 16'h3207; // 0x2e12
	13'h170a: q0 = 16'hd27c; // 0x2e14
	13'h170b: q0 = 16'h0080; // 0x2e16
	13'h170c: q0 = 16'h3081; // 0x2e18
	13'h170d: q0 = 16'h6018; // 0x2e1a
	13'h170e: q0 = 16'h0c55; // 0x2e1c
	13'h170f: q0 = 16'h0012; // 0x2e1e
	13'h1710: q0 = 16'h6f12; // 0x2e20
	13'h1711: q0 = 16'h0c55; // 0x2e22
	13'h1712: q0 = 16'h0036; // 0x2e24
	13'h1713: q0 = 16'h6e0c; // 0x2e26
	13'h1714: q0 = 16'h206d; // 0x2e28
	13'h1715: q0 = 16'h0022; // 0x2e2a
	13'h1716: q0 = 16'h3207; // 0x2e2c
	13'h1717: q0 = 16'hd27c; // 0x2e2e
	13'h1718: q0 = 16'hff80; // 0x2e30
	13'h1719: q0 = 16'h3081; // 0x2e32
	13'h171a: q0 = 16'h206d; // 0x2e34
	13'h171b: q0 = 16'h0022; // 0x2e36
	13'h171c: q0 = 16'h3146; // 0x2e38
	13'h171d: q0 = 16'h0002; // 0x2e3a
	13'h171e: q0 = 16'h082d; // 0x2e3c
	13'h171f: q0 = 16'h0002; // 0x2e3e
	13'h1720: q0 = 16'h000e; // 0x2e40
	13'h1721: q0 = 16'h661a; // 0x2e42
	13'h1722: q0 = 16'h0c55; // 0x2e44
	13'h1723: q0 = 16'h0012; // 0x2e46
	13'h1724: q0 = 16'h6f14; // 0x2e48
	13'h1725: q0 = 16'h0c55; // 0x2e4a
	13'h1726: q0 = 16'h0036; // 0x2e4c
	13'h1727: q0 = 16'h6e0e; // 0x2e4e
	13'h1728: q0 = 16'h206d; // 0x2e50
	13'h1729: q0 = 16'h0026; // 0x2e52
	13'h172a: q0 = 16'h3207; // 0x2e54
	13'h172b: q0 = 16'hd27c; // 0x2e56
	13'h172c: q0 = 16'hff80; // 0x2e58
	13'h172d: q0 = 16'h3081; // 0x2e5a
	13'h172e: q0 = 16'h6006; // 0x2e5c
	13'h172f: q0 = 16'h206d; // 0x2e5e
	13'h1730: q0 = 16'h0026; // 0x2e60
	13'h1731: q0 = 16'h3087; // 0x2e62
	13'h1732: q0 = 16'h206d; // 0x2e64
	13'h1733: q0 = 16'h0026; // 0x2e66
	13'h1734: q0 = 16'h3206; // 0x2e68
	13'h1735: q0 = 16'hd27c; // 0x2e6a
	13'h1736: q0 = 16'h0200; // 0x2e6c
	13'h1737: q0 = 16'h3141; // 0x2e6e
	13'h1738: q0 = 16'h0002; // 0x2e70
	13'h1739: q0 = 16'h4a9f; // 0x2e72
	13'h173a: q0 = 16'h4cdf; // 0x2e74
	13'h173b: q0 = 16'h20c0; // 0x2e76
	13'h173c: q0 = 16'h4e5e; // 0x2e78
	13'h173d: q0 = 16'h4e75; // 0x2e7a
	13'h173e: q0 = 16'h4e56; // 0x2e7c
	13'h173f: q0 = 16'h0000; // 0x2e7e
	13'h1740: q0 = 16'h48e7; // 0x2e80
	13'h1741: q0 = 16'h070c; // 0x2e82
	13'h1742: q0 = 16'h2c3c; // 0x2e84
	13'h1743: q0 = 16'h0000; // 0x2e86
	13'h1744: q0 = 16'h03e7; // 0x2e88
	13'h1745: q0 = 16'h2a7c; // 0x2e8a
	13'h1746: q0 = 16'h0001; // 0x2e8c
	13'h1747: q0 = 16'h89be; // 0x2e8e
	13'h1748: q0 = 16'h4247; // 0x2e90
	13'h1749: q0 = 16'hbe79; // 0x2e92
	13'h174a: q0 = 16'h0001; // 0x2e94
	13'h174b: q0 = 16'h7fbc; // 0x2e96
	13'h174c: q0 = 16'h6c18; // 0x2e98
	13'h174d: q0 = 16'h202d; // 0x2e9a
	13'h174e: q0 = 16'h002a; // 0x2e9c
	13'h174f: q0 = 16'hb086; // 0x2e9e
	13'h1750: q0 = 16'h6c06; // 0x2ea0
	13'h1751: q0 = 16'h2c2d; // 0x2ea2
	13'h1752: q0 = 16'h002a; // 0x2ea4
	13'h1753: q0 = 16'h284d; // 0x2ea6
	13'h1754: q0 = 16'hdbfc; // 0x2ea8
	13'h1755: q0 = 16'h0000; // 0x2eaa
	13'h1756: q0 = 16'h002e; // 0x2eac
	13'h1757: q0 = 16'h5247; // 0x2eae
	13'h1758: q0 = 16'h60e0; // 0x2eb0
	13'h1759: q0 = 16'h2a4c; // 0x2eb2
	13'h175a: q0 = 16'h42ad; // 0x2eb4
	13'h175b: q0 = 16'h002a; // 0x2eb6
	13'h175c: q0 = 16'h4a9f; // 0x2eb8
	13'h175d: q0 = 16'h4cdf; // 0x2eba
	13'h175e: q0 = 16'h30c0; // 0x2ebc
	13'h175f: q0 = 16'h4e5e; // 0x2ebe
	13'h1760: q0 = 16'h4e75; // 0x2ec0
	13'h1761: q0 = 16'h4e56; // 0x2ec2
	13'h1762: q0 = 16'hfffe; // 0x2ec4
	13'h1763: q0 = 16'h48e7; // 0x2ec6
	13'h1764: q0 = 16'h0104; // 0x2ec8
	13'h1765: q0 = 16'h2a6e; // 0x2eca
	13'h1766: q0 = 16'h0008; // 0x2ecc
	13'h1767: q0 = 16'h206d; // 0x2ece
	13'h1768: q0 = 16'h001e; // 0x2ed0
	13'h1769: q0 = 16'h317c; // 0x2ed2
	13'h176a: q0 = 16'h0030; // 0x2ed4
	13'h176b: q0 = 16'h0004; // 0x2ed6
	13'h176c: q0 = 16'h206d; // 0x2ed8
	13'h176d: q0 = 16'h0022; // 0x2eda
	13'h176e: q0 = 16'h317c; // 0x2edc
	13'h176f: q0 = 16'h0030; // 0x2ede
	13'h1770: q0 = 16'h0004; // 0x2ee0
	13'h1771: q0 = 16'h206d; // 0x2ee2
	13'h1772: q0 = 16'h0026; // 0x2ee4
	13'h1773: q0 = 16'h317c; // 0x2ee6
	13'h1774: q0 = 16'h0030; // 0x2ee8
	13'h1775: q0 = 16'h0004; // 0x2eea
	13'h1776: q0 = 16'h206d; // 0x2eec
	13'h1777: q0 = 16'h001e; // 0x2eee
	13'h1778: q0 = 16'h4250; // 0x2ef0
	13'h1779: q0 = 16'h206d; // 0x2ef2
	13'h177a: q0 = 16'h001e; // 0x2ef4
	13'h177b: q0 = 16'h4268; // 0x2ef6
	13'h177c: q0 = 16'h0002; // 0x2ef8
	13'h177d: q0 = 16'h206d; // 0x2efa
	13'h177e: q0 = 16'h001e; // 0x2efc
	13'h177f: q0 = 16'h4268; // 0x2efe
	13'h1780: q0 = 16'h0006; // 0x2f00
	13'h1781: q0 = 16'h206d; // 0x2f02
	13'h1782: q0 = 16'h0022; // 0x2f04
	13'h1783: q0 = 16'h4250; // 0x2f06
	13'h1784: q0 = 16'h206d; // 0x2f08
	13'h1785: q0 = 16'h0022; // 0x2f0a
	13'h1786: q0 = 16'h4268; // 0x2f0c
	13'h1787: q0 = 16'h0002; // 0x2f0e
	13'h1788: q0 = 16'h206d; // 0x2f10
	13'h1789: q0 = 16'h0022; // 0x2f12
	13'h178a: q0 = 16'h4268; // 0x2f14
	13'h178b: q0 = 16'h0006; // 0x2f16
	13'h178c: q0 = 16'h206d; // 0x2f18
	13'h178d: q0 = 16'h0026; // 0x2f1a
	13'h178e: q0 = 16'h4250; // 0x2f1c
	13'h178f: q0 = 16'h206d; // 0x2f1e
	13'h1790: q0 = 16'h0026; // 0x2f20
	13'h1791: q0 = 16'h4268; // 0x2f22
	13'h1792: q0 = 16'h0002; // 0x2f24
	13'h1793: q0 = 16'h206d; // 0x2f26
	13'h1794: q0 = 16'h0026; // 0x2f28
	13'h1795: q0 = 16'h4268; // 0x2f2a
	13'h1796: q0 = 16'h0006; // 0x2f2c
	13'h1797: q0 = 16'h4aad; // 0x2f2e
	13'h1798: q0 = 16'h0010; // 0x2f30
	13'h1799: q0 = 16'h670e; // 0x2f32
	13'h179a: q0 = 16'h2ead; // 0x2f34
	13'h179b: q0 = 16'h0010; // 0x2f36
	13'h179c: q0 = 16'h4eb9; // 0x2f38
	13'h179d: q0 = 16'h0000; // 0x2f3a
	13'h179e: q0 = 16'h3356; // 0x2f3c
	13'h179f: q0 = 16'h42ad; // 0x2f3e
	13'h17a0: q0 = 16'h0010; // 0x2f40
	13'h17a1: q0 = 16'h2079; // 0x2f42
	13'h17a2: q0 = 16'h0001; // 0x2f44
	13'h17a3: q0 = 16'h7fb8; // 0x2f46
	13'h17a4: q0 = 16'h3010; // 0x2f48
	13'h17a5: q0 = 16'heb40; // 0x2f4a
	13'h17a6: q0 = 16'h3d40; // 0x2f4c
	13'h17a7: q0 = 16'hfffe; // 0x2f4e
	13'h17a8: q0 = 16'h0c6e; // 0x2f50
	13'h17a9: q0 = 16'h00ff; // 0x2f52
	13'h17aa: q0 = 16'hfffe; // 0x2f54
	13'h17ab: q0 = 16'h6c12; // 0x2f56
	13'h17ac: q0 = 16'h303c; // 0x2f58
	13'h17ad: q0 = 16'h00ff; // 0x2f5a
	13'h17ae: q0 = 16'h906e; // 0x2f5c
	13'h17af: q0 = 16'hfffe; // 0x2f5e
	13'h17b0: q0 = 16'he240; // 0x2f60
	13'h17b1: q0 = 16'h48c0; // 0x2f62
	13'h17b2: q0 = 16'h2b40; // 0x2f64
	13'h17b3: q0 = 16'h002a; // 0x2f66
	13'h17b4: q0 = 16'h6004; // 0x2f68
	13'h17b5: q0 = 16'h42ad; // 0x2f6a
	13'h17b6: q0 = 16'h002a; // 0x2f6c
	13'h17b7: q0 = 16'h4a79; // 0x2f6e
	13'h17b8: q0 = 16'h0001; // 0x2f70
	13'h17b9: q0 = 16'h7faa; // 0x2f72
	13'h17ba: q0 = 16'h6708; // 0x2f74
	13'h17bb: q0 = 16'h2b7c; // 0x2f76
	13'h17bc: q0 = 16'h0000; // 0x2f78
	13'h17bd: q0 = 16'h2710; // 0x2f7a
	13'h17be: q0 = 16'h002a; // 0x2f7c
	13'h17bf: q0 = 16'h302d; // 0x2f7e
	13'h17c0: q0 = 16'h000e; // 0x2f80
	13'h17c1: q0 = 16'hc07c; // 0x2f82
	13'h17c2: q0 = 16'hf0f0; // 0x2f84
	13'h17c3: q0 = 16'h807c; // 0x2f86
	13'h17c4: q0 = 16'h0002; // 0x2f88
	13'h17c5: q0 = 16'h3b40; // 0x2f8a
	13'h17c6: q0 = 16'h000e; // 0x2f8c
	13'h17c7: q0 = 16'h5379; // 0x2f8e
	13'h17c8: q0 = 16'h0001; // 0x2f90
	13'h17c9: q0 = 16'h86d4; // 0x2f92
	13'h17ca: q0 = 16'h4a79; // 0x2f94
	13'h17cb: q0 = 16'h0001; // 0x2f96
	13'h17cc: q0 = 16'h86d4; // 0x2f98
	13'h17cd: q0 = 16'h660e; // 0x2f9a
	13'h17ce: q0 = 16'h4a79; // 0x2f9c
	13'h17cf: q0 = 16'h0001; // 0x2f9e
	13'h17d0: q0 = 16'h7faa; // 0x2fa0
	13'h17d1: q0 = 16'h6606; // 0x2fa2
	13'h17d2: q0 = 16'h4eb9; // 0x2fa4
	13'h17d3: q0 = 16'h0000; // 0x2fa6
	13'h17d4: q0 = 16'h2e7c; // 0x2fa8
	13'h17d5: q0 = 16'h4a9f; // 0x2faa
	13'h17d6: q0 = 16'h4cdf; // 0x2fac
	13'h17d7: q0 = 16'h2000; // 0x2fae
	13'h17d8: q0 = 16'h4e5e; // 0x2fb0
	13'h17d9: q0 = 16'h4e75; // 0x2fb2
	13'h17da: q0 = 16'h4e56; // 0x2fb4
	13'h17db: q0 = 16'hfffa; // 0x2fb6
	13'h17dc: q0 = 16'h48e7; // 0x2fb8
	13'h17dd: q0 = 16'h1f04; // 0x2fba
	13'h17de: q0 = 16'h4245; // 0x2fbc
	13'h17df: q0 = 16'h3e39; // 0x2fbe
	13'h17e0: q0 = 16'h0001; // 0x2fc0
	13'h17e1: q0 = 16'h86d6; // 0x2fc2
	13'h17e2: q0 = 16'h2a7c; // 0x2fc4
	13'h17e3: q0 = 16'h0001; // 0x2fc6
	13'h17e4: q0 = 16'h7bda; // 0x2fc8
	13'h17e5: q0 = 16'h4246; // 0x2fca
	13'h17e6: q0 = 16'hbc47; // 0x2fcc
	13'h17e7: q0 = 16'h6c00; // 0x2fce
	13'h17e8: q0 = 16'h0368; // 0x2fd0
	13'h17e9: q0 = 16'h4a6d; // 0x2fd2
	13'h17ea: q0 = 16'h0008; // 0x2fd4
	13'h17eb: q0 = 16'h6702; // 0x2fd6
	13'h17ec: q0 = 16'h5246; // 0x2fd8
	13'h17ed: q0 = 16'h0c6d; // 0x2fda
	13'h17ee: q0 = 16'h0003; // 0x2fdc
	13'h17ef: q0 = 16'h0008; // 0x2fde
	13'h17f0: q0 = 16'h6600; // 0x2fe0
	13'h17f1: q0 = 16'h022e; // 0x2fe2
	13'h17f2: q0 = 16'h4a6d; // 0x2fe4
	13'h17f3: q0 = 16'h0004; // 0x2fe6
	13'h17f4: q0 = 16'h6600; // 0x2fe8
	13'h17f5: q0 = 16'h01e0; // 0x2fea
	13'h17f6: q0 = 16'h4a79; // 0x2fec
	13'h17f7: q0 = 16'h0001; // 0x2fee
	13'h17f8: q0 = 16'h7bd6; // 0x2ff0
	13'h17f9: q0 = 16'h670c; // 0x2ff2
	13'h17fa: q0 = 16'h2e8d; // 0x2ff4
	13'h17fb: q0 = 16'h4eb9; // 0x2ff6
	13'h17fc: q0 = 16'h0000; // 0x2ff8
	13'h17fd: q0 = 16'h3356; // 0x2ffa
	13'h17fe: q0 = 16'h6000; // 0x2ffc
	13'h17ff: q0 = 16'h01c8; // 0x2ffe
	13'h1800: q0 = 16'h4a79; // 0x3000
	13'h1801: q0 = 16'h0001; // 0x3002
	13'h1802: q0 = 16'h7f2a; // 0x3004
	13'h1803: q0 = 16'h6700; // 0x3006
	13'h1804: q0 = 16'h00a0; // 0x3008
	13'h1805: q0 = 16'h3b7c; // 0x300a
	13'h1806: q0 = 16'h0005; // 0x300c
	13'h1807: q0 = 16'h0008; // 0x300e
	13'h1808: q0 = 16'h0c6d; // 0x3010
	13'h1809: q0 = 16'h0001; // 0x3012
	13'h180a: q0 = 16'h000a; // 0x3014
	13'h180b: q0 = 16'h6642; // 0x3016
	13'h180c: q0 = 16'h3806; // 0x3018
	13'h180d: q0 = 16'hc87c; // 0x301a
	13'h180e: q0 = 16'h0007; // 0x301c
	13'h180f: q0 = 16'h206d; // 0x301e
	13'h1810: q0 = 16'h0012; // 0x3020
	13'h1811: q0 = 16'h3204; // 0x3022
	13'h1812: q0 = 16'he341; // 0x3024
	13'h1813: q0 = 16'h48c1; // 0x3026
	13'h1814: q0 = 16'hd2bc; // 0x3028
	13'h1815: q0 = 16'h0000; // 0x302a
	13'h1816: q0 = 16'hc9a0; // 0x302c
	13'h1817: q0 = 16'h2241; // 0x302e
	13'h1818: q0 = 16'h3151; // 0x3030
	13'h1819: q0 = 16'h0004; // 0x3032
	13'h181a: q0 = 16'h206d; // 0x3034
	13'h181b: q0 = 16'h0012; // 0x3036
	13'h181c: q0 = 16'h226d; // 0x3038
	13'h181d: q0 = 16'h0012; // 0x303a
	13'h181e: q0 = 16'h3229; // 0x303c
	13'h181f: q0 = 16'h0006; // 0x303e
	13'h1820: q0 = 16'hc27c; // 0x3040
	13'h1821: q0 = 16'h003f; // 0x3042
	13'h1822: q0 = 16'h3404; // 0x3044
	13'h1823: q0 = 16'he342; // 0x3046
	13'h1824: q0 = 16'h48c2; // 0x3048
	13'h1825: q0 = 16'hd4bc; // 0x304a
	13'h1826: q0 = 16'h0000; // 0x304c
	13'h1827: q0 = 16'hc9b0; // 0x304e
	13'h1828: q0 = 16'h2442; // 0x3050
	13'h1829: q0 = 16'h8252; // 0x3052
	13'h182a: q0 = 16'h3141; // 0x3054
	13'h182b: q0 = 16'h0006; // 0x3056
	13'h182c: q0 = 16'h601a; // 0x3058
	13'h182d: q0 = 16'h206d; // 0x305a
	13'h182e: q0 = 16'h0012; // 0x305c
	13'h182f: q0 = 16'h226d; // 0x305e
	13'h1830: q0 = 16'h0016; // 0x3060
	13'h1831: q0 = 16'h3151; // 0x3062
	13'h1832: q0 = 16'h0004; // 0x3064
	13'h1833: q0 = 16'h206d; // 0x3066
	13'h1834: q0 = 16'h0012; // 0x3068
	13'h1835: q0 = 16'h226d; // 0x306a
	13'h1836: q0 = 16'h0016; // 0x306c
	13'h1837: q0 = 16'h3169; // 0x306e
	13'h1838: q0 = 16'h0002; // 0x3070
	13'h1839: q0 = 16'h0006; // 0x3072
	13'h183a: q0 = 16'h0c6d; // 0x3074
	13'h183b: q0 = 16'h0002; // 0x3076
	13'h183c: q0 = 16'h000a; // 0x3078
	13'h183d: q0 = 16'h6628; // 0x307a
	13'h183e: q0 = 16'h202d; // 0x307c
	13'h183f: q0 = 16'h0012; // 0x307e
	13'h1840: q0 = 16'h5c80; // 0x3080
	13'h1841: q0 = 16'h2e80; // 0x3082
	13'h1842: q0 = 16'h202d; // 0x3084
	13'h1843: q0 = 16'h0012; // 0x3086
	13'h1844: q0 = 16'h5880; // 0x3088
	13'h1845: q0 = 16'h2f00; // 0x308a
	13'h1846: q0 = 16'h3f2d; // 0x308c
	13'h1847: q0 = 16'h0002; // 0x308e
	13'h1848: q0 = 16'h3f15; // 0x3090
	13'h1849: q0 = 16'h4eb9; // 0x3092
	13'h184a: q0 = 16'h0000; // 0x3094
	13'h184b: q0 = 16'h0a1c; // 0x3096
	13'h184c: q0 = 16'h4a9f; // 0x3098
	13'h184d: q0 = 16'h3f00; // 0x309a
	13'h184e: q0 = 16'h4eb9; // 0x309c
	13'h184f: q0 = 16'h0000; // 0x309e
	13'h1850: q0 = 16'h3f1e; // 0x30a0
	13'h1851: q0 = 16'h5c4f; // 0x30a2
	13'h1852: q0 = 16'h6000; // 0x30a4
	13'h1853: q0 = 16'h0120; // 0x30a6
	13'h1854: q0 = 16'h206d; // 0x30a8
	13'h1855: q0 = 16'h0012; // 0x30aa
	13'h1856: q0 = 16'h3010; // 0x30ac
	13'h1857: q0 = 16'hd07c; // 0x30ae
	13'h1858: q0 = 16'h0200; // 0x30b0
	13'h1859: q0 = 16'h3d40; // 0x30b2
	13'h185a: q0 = 16'hfffc; // 0x30b4
	13'h185b: q0 = 16'h206d; // 0x30b6
	13'h185c: q0 = 16'h0012; // 0x30b8
	13'h185d: q0 = 16'h3028; // 0x30ba
	13'h185e: q0 = 16'h0002; // 0x30bc
	13'h185f: q0 = 16'hd07c; // 0x30be
	13'h1860: q0 = 16'h0200; // 0x30c0
	13'h1861: q0 = 16'h3d40; // 0x30c2
	13'h1862: q0 = 16'hfffa; // 0x30c4
	13'h1863: q0 = 16'h302e; // 0x30c6
	13'h1864: q0 = 16'hfffa; // 0x30c8
	13'h1865: q0 = 16'h4281; // 0x30ca
	13'h1866: q0 = 16'h720a; // 0x30cc
	13'h1867: q0 = 16'he260; // 0x30ce
	13'h1868: q0 = 16'heb40; // 0x30d0
	13'h1869: q0 = 16'h322e; // 0x30d2
	13'h186a: q0 = 16'hfffc; // 0x30d4
	13'h186b: q0 = 16'h4282; // 0x30d6
	13'h186c: q0 = 16'h740a; // 0x30d8
	13'h186d: q0 = 16'he461; // 0x30da
	13'h186e: q0 = 16'hd041; // 0x30dc
	13'h186f: q0 = 16'hd07c; // 0x30de
	13'h1870: q0 = 16'hfe00; // 0x30e0
	13'h1871: q0 = 16'h3d40; // 0x30e2
	13'h1872: q0 = 16'hfffe; // 0x30e4
	13'h1873: q0 = 16'h3ebc; // 0x30e6
	13'h1874: q0 = 16'h002c; // 0x30e8
	13'h1875: q0 = 16'h3f2e; // 0x30ea
	13'h1876: q0 = 16'hfffe; // 0x30ec
	13'h1877: q0 = 16'h3f2e; // 0x30ee
	13'h1878: q0 = 16'hfffa; // 0x30f0
	13'h1879: q0 = 16'h3f2e; // 0x30f2
	13'h187a: q0 = 16'hfffc; // 0x30f4
	13'h187b: q0 = 16'h4eb9; // 0x30f6
	13'h187c: q0 = 16'h0000; // 0x30f8
	13'h187d: q0 = 16'h3f80; // 0x30fa
	13'h187e: q0 = 16'h5c4f; // 0x30fc
	13'h187f: q0 = 16'h4a79; // 0x30fe
	13'h1880: q0 = 16'h0001; // 0x3100
	13'h1881: q0 = 16'h7f1c; // 0x3102
	13'h1882: q0 = 16'h6612; // 0x3104
	13'h1883: q0 = 16'h4a79; // 0x3106
	13'h1884: q0 = 16'h0001; // 0x3108
	13'h1885: q0 = 16'h7f1c; // 0x310a
	13'h1886: q0 = 16'h6616; // 0x310c
	13'h1887: q0 = 16'h0c79; // 0x310e
	13'h1888: q0 = 16'h000e; // 0x3110
	13'h1889: q0 = 16'h0001; // 0x3112
	13'h188a: q0 = 16'h7f1e; // 0x3114
	13'h188b: q0 = 16'h660c; // 0x3116
	13'h188c: q0 = 16'h2e8d; // 0x3118
	13'h188d: q0 = 16'h4eb9; // 0x311a
	13'h188e: q0 = 16'h0000; // 0x311c
	13'h188f: q0 = 16'h3356; // 0x311e
	13'h1890: q0 = 16'h6000; // 0x3120
	13'h1891: q0 = 16'h00a4; // 0x3122
	13'h1892: q0 = 16'h206d; // 0x3124
	13'h1893: q0 = 16'h0012; // 0x3126
	13'h1894: q0 = 16'h226d; // 0x3128
	13'h1895: q0 = 16'h0016; // 0x312a
	13'h1896: q0 = 16'h3151; // 0x312c
	13'h1897: q0 = 16'h0004; // 0x312e
	13'h1898: q0 = 16'h206d; // 0x3130
	13'h1899: q0 = 16'h0012; // 0x3132
	13'h189a: q0 = 16'h226d; // 0x3134
	13'h189b: q0 = 16'h0016; // 0x3136
	13'h189c: q0 = 16'h3169; // 0x3138
	13'h189d: q0 = 16'h0002; // 0x313a
	13'h189e: q0 = 16'h0006; // 0x313c
	13'h189f: q0 = 16'h3b7c; // 0x313e
	13'h18a0: q0 = 16'h0006; // 0x3140
	13'h18a1: q0 = 16'h0008; // 0x3142
	13'h18a2: q0 = 16'h0839; // 0x3144
	13'h18a3: q0 = 16'h0001; // 0x3146
	13'h18a4: q0 = 16'h0001; // 0x3148
	13'h18a5: q0 = 16'h7f1f; // 0x314a
	13'h18a6: q0 = 16'h6708; // 0x314c
	13'h18a7: q0 = 16'h3b7c; // 0x314e
	13'h18a8: q0 = 16'h0001; // 0x3150
	13'h18a9: q0 = 16'h001a; // 0x3152
	13'h18aa: q0 = 16'h6004; // 0x3154
	13'h18ab: q0 = 16'h426d; // 0x3156
	13'h18ac: q0 = 16'h001a; // 0x3158
	13'h18ad: q0 = 16'h3ebc; // 0x315a
	13'h18ae: q0 = 16'h0600; // 0x315c
	13'h18af: q0 = 16'h3f3c; // 0x315e
	13'h18b0: q0 = 16'h0200; // 0x3160
	13'h18b1: q0 = 16'h4eb9; // 0x3162
	13'h18b2: q0 = 16'h0000; // 0x3164
	13'h18b3: q0 = 16'h8e6c; // 0x3166
	13'h18b4: q0 = 16'h4a5f; // 0x3168
	13'h18b5: q0 = 16'h3a80; // 0x316a
	13'h18b6: q0 = 16'h0839; // 0x316c
	13'h18b7: q0 = 16'h0000; // 0x316e
	13'h18b8: q0 = 16'h0001; // 0x3170
	13'h18b9: q0 = 16'h7f1f; // 0x3172
	13'h18ba: q0 = 16'h6706; // 0x3174
	13'h18bb: q0 = 16'h3015; // 0x3176
	13'h18bc: q0 = 16'h4440; // 0x3178
	13'h18bd: q0 = 16'h3a80; // 0x317a
	13'h18be: q0 = 16'h426d; // 0x317c
	13'h18bf: q0 = 16'h0002; // 0x317e
	13'h18c0: q0 = 16'h0c6d; // 0x3180
	13'h18c1: q0 = 16'h0001; // 0x3182
	13'h18c2: q0 = 16'h000a; // 0x3184
	13'h18c3: q0 = 16'h6608; // 0x3186
	13'h18c4: q0 = 16'h3b7c; // 0x3188
	13'h18c5: q0 = 16'h7fff; // 0x318a
	13'h18c6: q0 = 16'h0004; // 0x318c
	13'h18c7: q0 = 16'h6030; // 0x318e
	13'h18c8: q0 = 16'h0c6d; // 0x3190
	13'h18c9: q0 = 16'h0002; // 0x3192
	13'h18ca: q0 = 16'h000a; // 0x3194
	13'h18cb: q0 = 16'h6628; // 0x3196
	13'h18cc: q0 = 16'h202d; // 0x3198
	13'h18cd: q0 = 16'h0012; // 0x319a
	13'h18ce: q0 = 16'h5c80; // 0x319c
	13'h18cf: q0 = 16'h2e80; // 0x319e
	13'h18d0: q0 = 16'h202d; // 0x31a0
	13'h18d1: q0 = 16'h0012; // 0x31a2
	13'h18d2: q0 = 16'h5880; // 0x31a4
	13'h18d3: q0 = 16'h2f00; // 0x31a6
	13'h18d4: q0 = 16'h3f2d; // 0x31a8
	13'h18d5: q0 = 16'h0002; // 0x31aa
	13'h18d6: q0 = 16'h3f15; // 0x31ac
	13'h18d7: q0 = 16'h4eb9; // 0x31ae
	13'h18d8: q0 = 16'h0000; // 0x31b0
	13'h18d9: q0 = 16'h0a1c; // 0x31b2
	13'h18da: q0 = 16'h4a9f; // 0x31b4
	13'h18db: q0 = 16'h3f00; // 0x31b6
	13'h18dc: q0 = 16'h4eb9; // 0x31b8
	13'h18dd: q0 = 16'h0000; // 0x31ba
	13'h18de: q0 = 16'h3f1e; // 0x31bc
	13'h18df: q0 = 16'h5c4f; // 0x31be
	13'h18e0: q0 = 16'h5279; // 0x31c0
	13'h18e1: q0 = 16'h0001; // 0x31c2
	13'h18e2: q0 = 16'h7f1e; // 0x31c4
	13'h18e3: q0 = 16'h6000; // 0x31c6
	13'h18e4: q0 = 16'h0166; // 0x31c8
	13'h18e5: q0 = 16'h0c6d; // 0x31ca
	13'h18e6: q0 = 16'h0003; // 0x31cc
	13'h18e7: q0 = 16'h000a; // 0x31ce
	13'h18e8: q0 = 16'h6620; // 0x31d0
	13'h18e9: q0 = 16'h0c6d; // 0x31d2
	13'h18ea: q0 = 16'h0004; // 0x31d4
	13'h18eb: q0 = 16'h0004; // 0x31d6
	13'h18ec: q0 = 16'h660e; // 0x31d8
	13'h18ed: q0 = 16'h206d; // 0x31da
	13'h18ee: q0 = 16'h0012; // 0x31dc
	13'h18ef: q0 = 16'h3179; // 0x31de
	13'h18f0: q0 = 16'h0000; // 0x31e0
	13'h18f1: q0 = 16'hc988; // 0x31e2
	13'h18f2: q0 = 16'h0004; // 0x31e4
	13'h18f3: q0 = 16'h6008; // 0x31e6
	13'h18f4: q0 = 16'h206d; // 0x31e8
	13'h18f5: q0 = 16'h0012; // 0x31ea
	13'h18f6: q0 = 16'h5268; // 0x31ec
	13'h18f7: q0 = 16'h0004; // 0x31ee
	13'h18f8: q0 = 16'h601a; // 0x31f0
	13'h18f9: q0 = 16'h206d; // 0x31f2
	13'h18fa: q0 = 16'h0012; // 0x31f4
	13'h18fb: q0 = 16'h322d; // 0x31f6
	13'h18fc: q0 = 16'h0004; // 0x31f8
	13'h18fd: q0 = 16'h5341; // 0x31fa
	13'h18fe: q0 = 16'he341; // 0x31fc
	13'h18ff: q0 = 16'h48c1; // 0x31fe
	13'h1900: q0 = 16'hd2bc; // 0x3200
	13'h1901: q0 = 16'h0000; // 0x3202
	13'h1902: q0 = 16'hc998; // 0x3204
	13'h1903: q0 = 16'h2241; // 0x3206
	13'h1904: q0 = 16'h3151; // 0x3208
	13'h1905: q0 = 16'h0004; // 0x320a
	13'h1906: q0 = 16'h536d; // 0x320c
	13'h1907: q0 = 16'h0004; // 0x320e
	13'h1908: q0 = 16'h0c6d; // 0x3210
	13'h1909: q0 = 16'h0002; // 0x3212
	13'h190a: q0 = 16'h0008; // 0x3214
	13'h190b: q0 = 16'h670a; // 0x3216
	13'h190c: q0 = 16'h0c6d; // 0x3218
	13'h190d: q0 = 16'h0006; // 0x321a
	13'h190e: q0 = 16'h0008; // 0x321c
	13'h190f: q0 = 16'h6600; // 0x321e
	13'h1910: q0 = 16'h010e; // 0x3220
	13'h1911: q0 = 16'h0c6d; // 0x3222
	13'h1912: q0 = 16'h0001; // 0x3224
	13'h1913: q0 = 16'h000a; // 0x3226
	13'h1914: q0 = 16'h6646; // 0x3228
	13'h1915: q0 = 16'h536d; // 0x322a
	13'h1916: q0 = 16'h0004; // 0x322c
	13'h1917: q0 = 16'h382d; // 0x322e
	13'h1918: q0 = 16'h0004; // 0x3230
	13'h1919: q0 = 16'hc87c; // 0x3232
	13'h191a: q0 = 16'h0007; // 0x3234
	13'h191b: q0 = 16'h206d; // 0x3236
	13'h191c: q0 = 16'h0012; // 0x3238
	13'h191d: q0 = 16'h3204; // 0x323a
	13'h191e: q0 = 16'he341; // 0x323c
	13'h191f: q0 = 16'h48c1; // 0x323e
	13'h1920: q0 = 16'hd2bc; // 0x3240
	13'h1921: q0 = 16'h0000; // 0x3242
	13'h1922: q0 = 16'hc9a0; // 0x3244
	13'h1923: q0 = 16'h2241; // 0x3246
	13'h1924: q0 = 16'h3151; // 0x3248
	13'h1925: q0 = 16'h0004; // 0x324a
	13'h1926: q0 = 16'h206d; // 0x324c
	13'h1927: q0 = 16'h0012; // 0x324e
	13'h1928: q0 = 16'h226d; // 0x3250
	13'h1929: q0 = 16'h0012; // 0x3252
	13'h192a: q0 = 16'h3229; // 0x3254
	13'h192b: q0 = 16'h0006; // 0x3256
	13'h192c: q0 = 16'hc27c; // 0x3258
	13'h192d: q0 = 16'h003f; // 0x325a
	13'h192e: q0 = 16'h3404; // 0x325c
	13'h192f: q0 = 16'he342; // 0x325e
	13'h1930: q0 = 16'h48c2; // 0x3260
	13'h1931: q0 = 16'hd4bc; // 0x3262
	13'h1932: q0 = 16'h0000; // 0x3264
	13'h1933: q0 = 16'hc9b0; // 0x3266
	13'h1934: q0 = 16'h2442; // 0x3268
	13'h1935: q0 = 16'h8252; // 0x326a
	13'h1936: q0 = 16'h3141; // 0x326c
	13'h1937: q0 = 16'h0006; // 0x326e
	13'h1938: q0 = 16'h3015; // 0x3270
	13'h1939: q0 = 16'h226d; // 0x3272
	13'h193a: q0 = 16'h0012; // 0x3274
	13'h193b: q0 = 16'hd151; // 0x3276
	13'h193c: q0 = 16'h0c6d; // 0x3278
	13'h193d: q0 = 16'h0006; // 0x327a
	13'h193e: q0 = 16'h0008; // 0x327c
	13'h193f: q0 = 16'h6700; // 0x327e
	13'h1940: q0 = 16'h00ae; // 0x3280
	13'h1941: q0 = 16'h206d; // 0x3282
	13'h1942: q0 = 16'h0012; // 0x3284
	13'h1943: q0 = 16'h3828; // 0x3286
	13'h1944: q0 = 16'h0002; // 0x3288
	13'h1945: q0 = 16'hd86d; // 0x328a
	13'h1946: q0 = 16'h0002; // 0x328c
	13'h1947: q0 = 16'h4a79; // 0x328e
	13'h1948: q0 = 16'h0001; // 0x3290
	13'h1949: q0 = 16'h7fc6; // 0x3292
	13'h194a: q0 = 16'h660a; // 0x3294
	13'h194b: q0 = 16'hb87c; // 0x3296
	13'h194c: q0 = 16'h7800; // 0x3298
	13'h194d: q0 = 16'h6f04; // 0x329a
	13'h194e: q0 = 16'h383c; // 0x329c
	13'h194f: q0 = 16'h7800; // 0x329e
	13'h1950: q0 = 16'h206d; // 0x32a0
	13'h1951: q0 = 16'h0012; // 0x32a2
	13'h1952: q0 = 16'h3144; // 0x32a4
	13'h1953: q0 = 16'h0002; // 0x32a6
	13'h1954: q0 = 16'h206d; // 0x32a8
	13'h1955: q0 = 16'h0012; // 0x32aa
	13'h1956: q0 = 16'h3010; // 0x32ac
	13'h1957: q0 = 16'hb06d; // 0x32ae
	13'h1958: q0 = 16'h001a; // 0x32b0
	13'h1959: q0 = 16'h6c0c; // 0x32b2
	13'h195a: q0 = 16'h302d; // 0x32b4
	13'h195b: q0 = 16'h001a; // 0x32b6
	13'h195c: q0 = 16'h226d; // 0x32b8
	13'h195d: q0 = 16'h0012; // 0x32ba
	13'h195e: q0 = 16'h9051; // 0x32bc
	13'h195f: q0 = 16'h600a; // 0x32be
	13'h1960: q0 = 16'h206d; // 0x32c0
	13'h1961: q0 = 16'h0012; // 0x32c2
	13'h1962: q0 = 16'h3010; // 0x32c4
	13'h1963: q0 = 16'h906d; // 0x32c6
	13'h1964: q0 = 16'h001a; // 0x32c8
	13'h1965: q0 = 16'hb06d; // 0x32ca
	13'h1966: q0 = 16'h0006; // 0x32cc
	13'h1967: q0 = 16'h6c5e; // 0x32ce
	13'h1968: q0 = 16'h206d; // 0x32d0
	13'h1969: q0 = 16'h0012; // 0x32d2
	13'h196a: q0 = 16'h3028; // 0x32d4
	13'h196b: q0 = 16'h0002; // 0x32d6
	13'h196c: q0 = 16'hb06d; // 0x32d8
	13'h196d: q0 = 16'h000c; // 0x32da
	13'h196e: q0 = 16'h6c0e; // 0x32dc
	13'h196f: q0 = 16'h302d; // 0x32de
	13'h1970: q0 = 16'h000c; // 0x32e0
	13'h1971: q0 = 16'h226d; // 0x32e2
	13'h1972: q0 = 16'h0012; // 0x32e4
	13'h1973: q0 = 16'h9069; // 0x32e6
	13'h1974: q0 = 16'h0002; // 0x32e8
	13'h1975: q0 = 16'h600c; // 0x32ea
	13'h1976: q0 = 16'h206d; // 0x32ec
	13'h1977: q0 = 16'h0012; // 0x32ee
	13'h1978: q0 = 16'h3028; // 0x32f0
	13'h1979: q0 = 16'h0002; // 0x32f2
	13'h197a: q0 = 16'h906d; // 0x32f4
	13'h197b: q0 = 16'h000c; // 0x32f6
	13'h197c: q0 = 16'hb06d; // 0x32f8
	13'h197d: q0 = 16'h0006; // 0x32fa
	13'h197e: q0 = 16'h6c30; // 0x32fc
	13'h197f: q0 = 16'h4a79; // 0x32fe
	13'h1980: q0 = 16'h0001; // 0x3300
	13'h1981: q0 = 16'h7fc6; // 0x3302
	13'h1982: q0 = 16'h6712; // 0x3304
	13'h1983: q0 = 16'h206d; // 0x3306
	13'h1984: q0 = 16'h0012; // 0x3308
	13'h1985: q0 = 16'h30ad; // 0x330a
	13'h1986: q0 = 16'h001a; // 0x330c
	13'h1987: q0 = 16'h206d; // 0x330e
	13'h1988: q0 = 16'h0012; // 0x3310
	13'h1989: q0 = 16'h316d; // 0x3312
	13'h198a: q0 = 16'h000c; // 0x3314
	13'h198b: q0 = 16'h0002; // 0x3316
	13'h198c: q0 = 16'h2e8d; // 0x3318
	13'h198d: q0 = 16'h4eb9; // 0x331a
	13'h198e: q0 = 16'h0000; // 0x331c
	13'h198f: q0 = 16'h3a1e; // 0x331e
	13'h1990: q0 = 16'h2ebc; // 0x3320
	13'h1991: q0 = 16'h0000; // 0x3322
	13'h1992: q0 = 16'hdfe6; // 0x3324
	13'h1993: q0 = 16'h4eb9; // 0x3326
	13'h1994: q0 = 16'h0000; // 0x3328
	13'h1995: q0 = 16'h7dd8; // 0x332a
	13'h1996: q0 = 16'h5245; // 0x332c
	13'h1997: q0 = 16'hdbfc; // 0x332e
	13'h1998: q0 = 16'h0000; // 0x3330
	13'h1999: q0 = 16'h001c; // 0x3332
	13'h199a: q0 = 16'h6000; // 0x3334
	13'h199b: q0 = 16'hfc96; // 0x3336
	13'h199c: q0 = 16'h4a79; // 0x3338
	13'h199d: q0 = 16'h0001; // 0x333a
	13'h199e: q0 = 16'h7bd6; // 0x333c
	13'h199f: q0 = 16'h670c; // 0x333e
	13'h19a0: q0 = 16'h4a45; // 0x3340
	13'h19a1: q0 = 16'h6f08; // 0x3342
	13'h19a2: q0 = 16'h3e85; // 0x3344
	13'h19a3: q0 = 16'h4eb9; // 0x3346
	13'h19a4: q0 = 16'h0000; // 0x3348
	13'h19a5: q0 = 16'h8ee8; // 0x334a
	13'h19a6: q0 = 16'h4a9f; // 0x334c
	13'h19a7: q0 = 16'h4cdf; // 0x334e
	13'h19a8: q0 = 16'h20f0; // 0x3350
	13'h19a9: q0 = 16'h4e5e; // 0x3352
	13'h19aa: q0 = 16'h4e75; // 0x3354
	13'h19ab: q0 = 16'h4e56; // 0x3356
	13'h19ac: q0 = 16'h0000; // 0x3358
	13'h19ad: q0 = 16'h48e7; // 0x335a
	13'h19ae: q0 = 16'h0104; // 0x335c
	13'h19af: q0 = 16'h2a6e; // 0x335e
	13'h19b0: q0 = 16'h0008; // 0x3360
	13'h19b1: q0 = 16'h426d; // 0x3362
	13'h19b2: q0 = 16'h0008; // 0x3364
	13'h19b3: q0 = 16'h206d; // 0x3366
	13'h19b4: q0 = 16'h0012; // 0x3368
	13'h19b5: q0 = 16'h317c; // 0x336a
	13'h19b6: q0 = 16'h0030; // 0x336c
	13'h19b7: q0 = 16'h0004; // 0x336e
	13'h19b8: q0 = 16'h206d; // 0x3370
	13'h19b9: q0 = 16'h0012; // 0x3372
	13'h19ba: q0 = 16'h4250; // 0x3374
	13'h19bb: q0 = 16'h206d; // 0x3376
	13'h19bc: q0 = 16'h0012; // 0x3378
	13'h19bd: q0 = 16'h4268; // 0x337a
	13'h19be: q0 = 16'h0002; // 0x337c
	13'h19bf: q0 = 16'h206d; // 0x337e
	13'h19c0: q0 = 16'h0012; // 0x3380
	13'h19c1: q0 = 16'h4268; // 0x3382
	13'h19c2: q0 = 16'h0006; // 0x3384
	13'h19c3: q0 = 16'h5379; // 0x3386
	13'h19c4: q0 = 16'h0001; // 0x3388
	13'h19c5: q0 = 16'h86d6; // 0x338a
	13'h19c6: q0 = 16'h4a9f; // 0x338c
	13'h19c7: q0 = 16'h4cdf; // 0x338e
	13'h19c8: q0 = 16'h2000; // 0x3390
	13'h19c9: q0 = 16'h4e5e; // 0x3392
	13'h19ca: q0 = 16'h4e75; // 0x3394
	13'h19cb: q0 = 16'h4e56; // 0x3396
	13'h19cc: q0 = 16'h0000; // 0x3398
	13'h19cd: q0 = 16'h48e7; // 0x339a
	13'h19ce: q0 = 16'h0304; // 0x339c
	13'h19cf: q0 = 16'h2a7c; // 0x339e
	13'h19d0: q0 = 16'h0001; // 0x33a0
	13'h19d1: q0 = 16'h7bda; // 0x33a2
	13'h19d2: q0 = 16'h4247; // 0x33a4
	13'h19d3: q0 = 16'hbe79; // 0x33a6
	13'h19d4: q0 = 16'h0001; // 0x33a8
	13'h19d5: q0 = 16'h86d6; // 0x33aa
	13'h19d6: q0 = 16'h6c2c; // 0x33ac
	13'h19d7: q0 = 16'h4a6d; // 0x33ae
	13'h19d8: q0 = 16'h0008; // 0x33b0
	13'h19d9: q0 = 16'h671e; // 0x33b2
	13'h19da: q0 = 16'h0c6d; // 0x33b4
	13'h19db: q0 = 16'h0002; // 0x33b6
	13'h19dc: q0 = 16'h0008; // 0x33b8
	13'h19dd: q0 = 16'h6710; // 0x33ba
	13'h19de: q0 = 16'h0c6d; // 0x33bc
	13'h19df: q0 = 16'h0003; // 0x33be
	13'h19e0: q0 = 16'h0008; // 0x33c0
	13'h19e1: q0 = 16'h6708; // 0x33c2
	13'h19e2: q0 = 16'h0c6d; // 0x33c4
	13'h19e3: q0 = 16'h0004; // 0x33c6
	13'h19e4: q0 = 16'h0008; // 0x33c8
	13'h19e5: q0 = 16'h6604; // 0x33ca
	13'h19e6: q0 = 16'h4240; // 0x33cc
	13'h19e7: q0 = 16'h600c; // 0x33ce
	13'h19e8: q0 = 16'h5247; // 0x33d0
	13'h19e9: q0 = 16'hdbfc; // 0x33d2
	13'h19ea: q0 = 16'h0000; // 0x33d4
	13'h19eb: q0 = 16'h001c; // 0x33d6
	13'h19ec: q0 = 16'h60cc; // 0x33d8
	13'h19ed: q0 = 16'h7001; // 0x33da
	13'h19ee: q0 = 16'h4a9f; // 0x33dc
	13'h19ef: q0 = 16'h4cdf; // 0x33de
	13'h19f0: q0 = 16'h2080; // 0x33e0
	13'h19f1: q0 = 16'h4e5e; // 0x33e2
	13'h19f2: q0 = 16'h4e75; // 0x33e4
	13'h19f3: q0 = 16'h4e56; // 0x33e6
	13'h19f4: q0 = 16'h0000; // 0x33e8
	13'h19f5: q0 = 16'h48e7; // 0x33ea
	13'h19f6: q0 = 16'h0304; // 0x33ec
	13'h19f7: q0 = 16'h2a7c; // 0x33ee
	13'h19f8: q0 = 16'h0001; // 0x33f0
	13'h19f9: q0 = 16'h7bda; // 0x33f2
	13'h19fa: q0 = 16'h4247; // 0x33f4
	13'h19fb: q0 = 16'hbe7c; // 0x33f6
	13'h19fc: q0 = 16'h001a; // 0x33f8
	13'h19fd: q0 = 16'h6c2e; // 0x33fa
	13'h19fe: q0 = 16'h206d; // 0x33fc
	13'h19ff: q0 = 16'h0012; // 0x33fe
	13'h1a00: q0 = 16'h4250; // 0x3400
	13'h1a01: q0 = 16'h206d; // 0x3402
	13'h1a02: q0 = 16'h0012; // 0x3404
	13'h1a03: q0 = 16'h4268; // 0x3406
	13'h1a04: q0 = 16'h0002; // 0x3408
	13'h1a05: q0 = 16'h206d; // 0x340a
	13'h1a06: q0 = 16'h0012; // 0x340c
	13'h1a07: q0 = 16'h317c; // 0x340e
	13'h1a08: q0 = 16'h0030; // 0x3410
	13'h1a09: q0 = 16'h0004; // 0x3412
	13'h1a0a: q0 = 16'h206d; // 0x3414
	13'h1a0b: q0 = 16'h0012; // 0x3416
	13'h1a0c: q0 = 16'h4268; // 0x3418
	13'h1a0d: q0 = 16'h0006; // 0x341a
	13'h1a0e: q0 = 16'h426d; // 0x341c
	13'h1a0f: q0 = 16'h0008; // 0x341e
	13'h1a10: q0 = 16'hdbfc; // 0x3420
	13'h1a11: q0 = 16'h0000; // 0x3422
	13'h1a12: q0 = 16'h001c; // 0x3424
	13'h1a13: q0 = 16'h5247; // 0x3426
	13'h1a14: q0 = 16'h60cc; // 0x3428
	13'h1a15: q0 = 16'h4a9f; // 0x342a
	13'h1a16: q0 = 16'h4cdf; // 0x342c
	13'h1a17: q0 = 16'h2080; // 0x342e
	13'h1a18: q0 = 16'h4e5e; // 0x3430
	13'h1a19: q0 = 16'h4e75; // 0x3432
	13'h1a1a: q0 = 16'h4e56; // 0x3434
	13'h1a1b: q0 = 16'h0000; // 0x3436
	13'h1a1c: q0 = 16'h48e7; // 0x3438
	13'h1a1d: q0 = 16'h1f04; // 0x343a
	13'h1a1e: q0 = 16'h3e39; // 0x343c
	13'h1a1f: q0 = 16'h0001; // 0x343e
	13'h1a20: q0 = 16'h86d6; // 0x3440
	13'h1a21: q0 = 16'h0c79; // 0x3442
	13'h1a22: q0 = 16'h0001; // 0x3444
	13'h1a23: q0 = 16'h0001; // 0x3446
	13'h1a24: q0 = 16'h757c; // 0x3448
	13'h1a25: q0 = 16'h6f06; // 0x344a
	13'h1a26: q0 = 16'h54b9; // 0x344c
	13'h1a27: q0 = 16'h0001; // 0x344e
	13'h1a28: q0 = 16'h7eb2; // 0x3450
	13'h1a29: q0 = 16'h2a7c; // 0x3452
	13'h1a2a: q0 = 16'h0001; // 0x3454
	13'h1a2b: q0 = 16'h7bda; // 0x3456
	13'h1a2c: q0 = 16'h4246; // 0x3458
	13'h1a2d: q0 = 16'hbc47; // 0x345a
	13'h1a2e: q0 = 16'h6c00; // 0x345c
	13'h1a2f: q0 = 16'h0270; // 0x345e
	13'h1a30: q0 = 16'h4a6d; // 0x3460
	13'h1a31: q0 = 16'h0008; // 0x3462
	13'h1a32: q0 = 16'h6702; // 0x3464
	13'h1a33: q0 = 16'h5246; // 0x3466
	13'h1a34: q0 = 16'h0c6d; // 0x3468
	13'h1a35: q0 = 16'h0003; // 0x346a
	13'h1a36: q0 = 16'h0008; // 0x346c
	13'h1a37: q0 = 16'h6600; // 0x346e
	13'h1a38: q0 = 16'h00ae; // 0x3470
	13'h1a39: q0 = 16'h4a6d; // 0x3472
	13'h1a3a: q0 = 16'h0004; // 0x3474
	13'h1a3b: q0 = 16'h665c; // 0x3476
	13'h1a3c: q0 = 16'h4aad; // 0x3478
	13'h1a3d: q0 = 16'h000e; // 0x347a
	13'h1a3e: q0 = 16'h664e; // 0x347c
	13'h1a3f: q0 = 16'h4a79; // 0x347e
	13'h1a40: q0 = 16'h0001; // 0x3480
	13'h1a41: q0 = 16'h7f20; // 0x3482
	13'h1a42: q0 = 16'h6646; // 0x3484
	13'h1a43: q0 = 16'h0c79; // 0x3486
	13'h1a44: q0 = 16'h000a; // 0x3488
	13'h1a45: q0 = 16'h0001; // 0x348a
	13'h1a46: q0 = 16'h7ba0; // 0x348c
	13'h1a47: q0 = 16'h6c06; // 0x348e
	13'h1a48: q0 = 16'h5279; // 0x3490
	13'h1a49: q0 = 16'h0001; // 0x3492
	13'h1a4a: q0 = 16'h7ba0; // 0x3494
	13'h1a4b: q0 = 16'h3eb9; // 0x3496
	13'h1a4c: q0 = 16'h0001; // 0x3498
	13'h1a4d: q0 = 16'h7ba0; // 0x349a
	13'h1a4e: q0 = 16'h4eb9; // 0x349c
	13'h1a4f: q0 = 16'h0000; // 0x349e
	13'h1a50: q0 = 16'h8ee8; // 0x34a0
	13'h1a51: q0 = 16'h206d; // 0x34a2
	13'h1a52: q0 = 16'h0012; // 0x34a4
	13'h1a53: q0 = 16'h3239; // 0x34a6
	13'h1a54: q0 = 16'h0001; // 0x34a8
	13'h1a55: q0 = 16'h7ba0; // 0x34aa
	13'h1a56: q0 = 16'hd27c; // 0x34ac
	13'h1a57: q0 = 16'h0042; // 0x34ae
	13'h1a58: q0 = 16'h3141; // 0x34b0
	13'h1a59: q0 = 16'h0004; // 0x34b2
	13'h1a5a: q0 = 16'h206d; // 0x34b4
	13'h1a5b: q0 = 16'h0012; // 0x34b6
	13'h1a5c: q0 = 16'h317c; // 0x34b8
	13'h1a5d: q0 = 16'h001f; // 0x34ba
	13'h1a5e: q0 = 16'h0006; // 0x34bc
	13'h1a5f: q0 = 16'h3b7c; // 0x34be
	13'h1a60: q0 = 16'h0004; // 0x34c0
	13'h1a61: q0 = 16'h0008; // 0x34c2
	13'h1a62: q0 = 16'h3b7c; // 0x34c4
	13'h1a63: q0 = 16'h000a; // 0x34c6
	13'h1a64: q0 = 16'h0004; // 0x34c8
	13'h1a65: q0 = 16'h6004; // 0x34ca
	13'h1a66: q0 = 16'h6000; // 0x34cc
	13'h1a67: q0 = 16'h01ee; // 0x34ce
	13'h1a68: q0 = 16'h6000; // 0x34d0
	13'h1a69: q0 = 16'h01f2; // 0x34d2
	13'h1a6a: q0 = 16'h0c6d; // 0x34d4
	13'h1a6b: q0 = 16'h0003; // 0x34d6
	13'h1a6c: q0 = 16'h000a; // 0x34d8
	13'h1a6d: q0 = 16'h6620; // 0x34da
	13'h1a6e: q0 = 16'h0c6d; // 0x34dc
	13'h1a6f: q0 = 16'h0004; // 0x34de
	13'h1a70: q0 = 16'h0004; // 0x34e0
	13'h1a71: q0 = 16'h660e; // 0x34e2
	13'h1a72: q0 = 16'h206d; // 0x34e4
	13'h1a73: q0 = 16'h0012; // 0x34e6
	13'h1a74: q0 = 16'h3179; // 0x34e8
	13'h1a75: q0 = 16'h0000; // 0x34ea
	13'h1a76: q0 = 16'hc988; // 0x34ec
	13'h1a77: q0 = 16'h0004; // 0x34ee
	13'h1a78: q0 = 16'h6008; // 0x34f0
	13'h1a79: q0 = 16'h206d; // 0x34f2
	13'h1a7a: q0 = 16'h0012; // 0x34f4
	13'h1a7b: q0 = 16'h5268; // 0x34f6
	13'h1a7c: q0 = 16'h0004; // 0x34f8
	13'h1a7d: q0 = 16'h601a; // 0x34fa
	13'h1a7e: q0 = 16'h206d; // 0x34fc
	13'h1a7f: q0 = 16'h0012; // 0x34fe
	13'h1a80: q0 = 16'h322d; // 0x3500
	13'h1a81: q0 = 16'h0004; // 0x3502
	13'h1a82: q0 = 16'h5341; // 0x3504
	13'h1a83: q0 = 16'he341; // 0x3506
	13'h1a84: q0 = 16'h48c1; // 0x3508
	13'h1a85: q0 = 16'hd2bc; // 0x350a
	13'h1a86: q0 = 16'h0000; // 0x350c
	13'h1a87: q0 = 16'hc998; // 0x350e
	13'h1a88: q0 = 16'h2241; // 0x3510
	13'h1a89: q0 = 16'h3151; // 0x3512
	13'h1a8a: q0 = 16'h0004; // 0x3514
	13'h1a8b: q0 = 16'h536d; // 0x3516
	13'h1a8c: q0 = 16'h0004; // 0x3518
	13'h1a8d: q0 = 16'h6000; // 0x351a
	13'h1a8e: q0 = 16'h00f0; // 0x351c
	13'h1a8f: q0 = 16'h0c6d; // 0x351e
	13'h1a90: q0 = 16'h0004; // 0x3520
	13'h1a91: q0 = 16'h0008; // 0x3522
	13'h1a92: q0 = 16'h6614; // 0x3524
	13'h1a93: q0 = 16'h4a6d; // 0x3526
	13'h1a94: q0 = 16'h0004; // 0x3528
	13'h1a95: q0 = 16'h6700; // 0x352a
	13'h1a96: q0 = 16'h0190; // 0x352c
	13'h1a97: q0 = 16'h536d; // 0x352e
	13'h1a98: q0 = 16'h0004; // 0x3530
	13'h1a99: q0 = 16'h6000; // 0x3532
	13'h1a9a: q0 = 16'h0190; // 0x3534
	13'h1a9b: q0 = 16'h6000; // 0x3536
	13'h1a9c: q0 = 16'h00d4; // 0x3538
	13'h1a9d: q0 = 16'h0c6d; // 0x353a
	13'h1a9e: q0 = 16'h0002; // 0x353c
	13'h1a9f: q0 = 16'h0008; // 0x353e
	13'h1aa0: q0 = 16'h670a; // 0x3540
	13'h1aa1: q0 = 16'h0c6d; // 0x3542
	13'h1aa2: q0 = 16'h0006; // 0x3544
	13'h1aa3: q0 = 16'h0008; // 0x3546
	13'h1aa4: q0 = 16'h6600; // 0x3548
	13'h1aa5: q0 = 16'h00be; // 0x354a
	13'h1aa6: q0 = 16'h0c6d; // 0x354c
	13'h1aa7: q0 = 16'h0002; // 0x354e
	13'h1aa8: q0 = 16'h0008; // 0x3550
	13'h1aa9: q0 = 16'h6608; // 0x3552
	13'h1aaa: q0 = 16'h4a6d; // 0x3554
	13'h1aab: q0 = 16'h0004; // 0x3556
	13'h1aac: q0 = 16'h6700; // 0x3558
	13'h1aad: q0 = 16'h0162; // 0x355a
	13'h1aae: q0 = 16'h0c6d; // 0x355c
	13'h1aaf: q0 = 16'h0006; // 0x355e
	13'h1ab0: q0 = 16'h0008; // 0x3560
	13'h1ab1: q0 = 16'h6608; // 0x3562
	13'h1ab2: q0 = 16'h3015; // 0x3564
	13'h1ab3: q0 = 16'h226d; // 0x3566
	13'h1ab4: q0 = 16'h0012; // 0x3568
	13'h1ab5: q0 = 16'hd151; // 0x356a
	13'h1ab6: q0 = 16'h536d; // 0x356c
	13'h1ab7: q0 = 16'h0004; // 0x356e
	13'h1ab8: q0 = 16'h0c6d; // 0x3570
	13'h1ab9: q0 = 16'h0001; // 0x3572
	13'h1aba: q0 = 16'h000a; // 0x3574
	13'h1abb: q0 = 16'h6642; // 0x3576
	13'h1abc: q0 = 16'h382d; // 0x3578
	13'h1abd: q0 = 16'h0004; // 0x357a
	13'h1abe: q0 = 16'hc87c; // 0x357c
	13'h1abf: q0 = 16'h0007; // 0x357e
	13'h1ac0: q0 = 16'h206d; // 0x3580
	13'h1ac1: q0 = 16'h0012; // 0x3582
	13'h1ac2: q0 = 16'h3204; // 0x3584
	13'h1ac3: q0 = 16'he341; // 0x3586
	13'h1ac4: q0 = 16'h48c1; // 0x3588
	13'h1ac5: q0 = 16'hd2bc; // 0x358a
	13'h1ac6: q0 = 16'h0000; // 0x358c
	13'h1ac7: q0 = 16'hc9a0; // 0x358e
	13'h1ac8: q0 = 16'h2241; // 0x3590
	13'h1ac9: q0 = 16'h3151; // 0x3592
	13'h1aca: q0 = 16'h0004; // 0x3594
	13'h1acb: q0 = 16'h206d; // 0x3596
	13'h1acc: q0 = 16'h0012; // 0x3598
	13'h1acd: q0 = 16'h226d; // 0x359a
	13'h1ace: q0 = 16'h0012; // 0x359c
	13'h1acf: q0 = 16'h3229; // 0x359e
	13'h1ad0: q0 = 16'h0006; // 0x35a0
	13'h1ad1: q0 = 16'hc27c; // 0x35a2
	13'h1ad2: q0 = 16'h003f; // 0x35a4
	13'h1ad3: q0 = 16'h3404; // 0x35a6
	13'h1ad4: q0 = 16'he342; // 0x35a8
	13'h1ad5: q0 = 16'h48c2; // 0x35aa
	13'h1ad6: q0 = 16'hd4bc; // 0x35ac
	13'h1ad7: q0 = 16'h0000; // 0x35ae
	13'h1ad8: q0 = 16'hc9b0; // 0x35b0
	13'h1ad9: q0 = 16'h2442; // 0x35b2
	13'h1ada: q0 = 16'h8252; // 0x35b4
	13'h1adb: q0 = 16'h3141; // 0x35b6
	13'h1adc: q0 = 16'h0006; // 0x35b8
	13'h1add: q0 = 16'h0c6d; // 0x35ba
	13'h1ade: q0 = 16'h0006; // 0x35bc
	13'h1adf: q0 = 16'h0008; // 0x35be
	13'h1ae0: q0 = 16'h6700; // 0x35c0
	13'h1ae1: q0 = 16'h0102; // 0x35c2
	13'h1ae2: q0 = 16'h0c6d; // 0x35c4
	13'h1ae3: q0 = 16'h0002; // 0x35c6
	13'h1ae4: q0 = 16'h0008; // 0x35c8
	13'h1ae5: q0 = 16'h663a; // 0x35ca
	13'h1ae6: q0 = 16'h0c6d; // 0x35cc
	13'h1ae7: q0 = 16'h0003; // 0x35ce
	13'h1ae8: q0 = 16'h000a; // 0x35d0
	13'h1ae9: q0 = 16'h6632; // 0x35d2
	13'h1aea: q0 = 16'h382d; // 0x35d4
	13'h1aeb: q0 = 16'h0004; // 0x35d6
	13'h1aec: q0 = 16'he444; // 0x35d8
	13'h1aed: q0 = 16'h206d; // 0x35da
	13'h1aee: q0 = 16'h0012; // 0x35dc
	13'h1aef: q0 = 16'h7203; // 0x35de
	13'h1af0: q0 = 16'h9244; // 0x35e0
	13'h1af1: q0 = 16'he341; // 0x35e2
	13'h1af2: q0 = 16'h48c1; // 0x35e4
	13'h1af3: q0 = 16'hd2bc; // 0x35e6
	13'h1af4: q0 = 16'h0000; // 0x35e8
	13'h1af5: q0 = 16'hc988; // 0x35ea
	13'h1af6: q0 = 16'h2241; // 0x35ec
	13'h1af7: q0 = 16'h3151; // 0x35ee
	13'h1af8: q0 = 16'h0004; // 0x35f0
	13'h1af9: q0 = 16'h7003; // 0x35f2
	13'h1afa: q0 = 16'h9044; // 0x35f4
	13'h1afb: q0 = 16'he340; // 0x35f6
	13'h1afc: q0 = 16'h48c0; // 0x35f8
	13'h1afd: q0 = 16'hd0bc; // 0x35fa
	13'h1afe: q0 = 16'h0000; // 0x35fc
	13'h1aff: q0 = 16'hc990; // 0x35fe
	13'h1b00: q0 = 16'h2040; // 0x3600
	13'h1b01: q0 = 16'h3b50; // 0x3602
	13'h1b02: q0 = 16'h0006; // 0x3604
	13'h1b03: q0 = 16'h6004; // 0x3606
	13'h1b04: q0 = 16'h6000; // 0x3608
	13'h1b05: q0 = 16'h00ba; // 0x360a
	13'h1b06: q0 = 16'h206d; // 0x360c
	13'h1b07: q0 = 16'h0012; // 0x360e
	13'h1b08: q0 = 16'h3a10; // 0x3610
	13'h1b09: q0 = 16'hda55; // 0x3612
	13'h1b0a: q0 = 16'hba7c; // 0x3614
	13'h1b0b: q0 = 16'h0080; // 0x3616
	13'h1b0c: q0 = 16'h6c10; // 0x3618
	13'h1b0d: q0 = 16'h4a55; // 0x361a
	13'h1b0e: q0 = 16'h6f06; // 0x361c
	13'h1b0f: q0 = 16'h3a3c; // 0x361e
	13'h1b10: q0 = 16'h0080; // 0x3620
	13'h1b11: q0 = 16'h6004; // 0x3622
	13'h1b12: q0 = 16'h6000; // 0x3624
	13'h1b13: q0 = 16'h0096; // 0x3626
	13'h1b14: q0 = 16'h6014; // 0x3628
	13'h1b15: q0 = 16'hba7c; // 0x362a
	13'h1b16: q0 = 16'h7880; // 0x362c
	13'h1b17: q0 = 16'h6f0e; // 0x362e
	13'h1b18: q0 = 16'h4a55; // 0x3630
	13'h1b19: q0 = 16'h6c06; // 0x3632
	13'h1b1a: q0 = 16'h3a3c; // 0x3634
	13'h1b1b: q0 = 16'h7880; // 0x3636
	13'h1b1c: q0 = 16'h6004; // 0x3638
	13'h1b1d: q0 = 16'h6000; // 0x363a
	13'h1b1e: q0 = 16'h0080; // 0x363c
	13'h1b1f: q0 = 16'h206d; // 0x363e
	13'h1b20: q0 = 16'h0012; // 0x3640
	13'h1b21: q0 = 16'h3085; // 0x3642
	13'h1b22: q0 = 16'h206d; // 0x3644
	13'h1b23: q0 = 16'h0012; // 0x3646
	13'h1b24: q0 = 16'h3a28; // 0x3648
	13'h1b25: q0 = 16'h0002; // 0x364a
	13'h1b26: q0 = 16'hda6d; // 0x364c
	13'h1b27: q0 = 16'h0002; // 0x364e
	13'h1b28: q0 = 16'hba7c; // 0x3650
	13'h1b29: q0 = 16'h1280; // 0x3652
	13'h1b2a: q0 = 16'h6d66; // 0x3654
	13'h1b2b: q0 = 16'hba7c; // 0x3656
	13'h1b2c: q0 = 16'h7800; // 0x3658
	13'h1b2d: q0 = 16'h6e60; // 0x365a
	13'h1b2e: q0 = 16'h206d; // 0x365c
	13'h1b2f: q0 = 16'h0012; // 0x365e
	13'h1b30: q0 = 16'h3145; // 0x3660
	13'h1b31: q0 = 16'h0002; // 0x3662
	13'h1b32: q0 = 16'h4eb9; // 0x3664
	13'h1b33: q0 = 16'h0000; // 0x3666
	13'h1b34: q0 = 16'h4ec6; // 0x3668
	13'h1b35: q0 = 16'hb07c; // 0x366a
	13'h1b36: q0 = 16'h0002; // 0x366c
	13'h1b37: q0 = 16'h664a; // 0x366e
	13'h1b38: q0 = 16'h2039; // 0x3670
	13'h1b39: q0 = 16'h0000; // 0x3672
	13'h1b3a: q0 = 16'hc8d2; // 0x3674
	13'h1b3b: q0 = 16'he380; // 0x3676
	13'h1b3c: q0 = 16'hb0ad; // 0x3678
	13'h1b3d: q0 = 16'h000e; // 0x367a
	13'h1b3e: q0 = 16'h663c; // 0x367c
	13'h1b3f: q0 = 16'h4eb9; // 0x367e
	13'h1b40: q0 = 16'h0000; // 0x3680
	13'h1b41: q0 = 16'h4ee2; // 0x3682
	13'h1b42: q0 = 16'h3e80; // 0x3684
	13'h1b43: q0 = 16'h206d; // 0x3686
	13'h1b44: q0 = 16'h0012; // 0x3688
	13'h1b45: q0 = 16'h3010; // 0x368a
	13'h1b46: q0 = 16'h9157; // 0x368c
	13'h1b47: q0 = 16'h4eb9; // 0x368e
	13'h1b48: q0 = 16'h0000; // 0x3690
	13'h1b49: q0 = 16'h09a2; // 0x3692
	13'h1b4a: q0 = 16'hb07c; // 0x3694
	13'h1b4b: q0 = 16'h0480; // 0x3696
	13'h1b4c: q0 = 16'h6c2a; // 0x3698
	13'h1b4d: q0 = 16'h4eb9; // 0x369a
	13'h1b4e: q0 = 16'h0000; // 0x369c
	13'h1b4f: q0 = 16'h4f30; // 0x369e
	13'h1b50: q0 = 16'h3e80; // 0x36a0
	13'h1b51: q0 = 16'h206d; // 0x36a2
	13'h1b52: q0 = 16'h0012; // 0x36a4
	13'h1b53: q0 = 16'h3028; // 0x36a6
	13'h1b54: q0 = 16'h0002; // 0x36a8
	13'h1b55: q0 = 16'h9157; // 0x36aa
	13'h1b56: q0 = 16'h4eb9; // 0x36ac
	13'h1b57: q0 = 16'h0000; // 0x36ae
	13'h1b58: q0 = 16'h09a2; // 0x36b0
	13'h1b59: q0 = 16'hb07c; // 0x36b2
	13'h1b5a: q0 = 16'h0480; // 0x36b4
	13'h1b5b: q0 = 16'h6c0c; // 0x36b6
	13'h1b5c: q0 = 16'h6002; // 0x36b8
	13'h1b5d: q0 = 16'h6008; // 0x36ba
	13'h1b5e: q0 = 16'h2e8d; // 0x36bc
	13'h1b5f: q0 = 16'h4eb9; // 0x36be
	13'h1b60: q0 = 16'h0000; // 0x36c0
	13'h1b61: q0 = 16'h3356; // 0x36c2
	13'h1b62: q0 = 16'hdbfc; // 0x36c4
	13'h1b63: q0 = 16'h0000; // 0x36c6
	13'h1b64: q0 = 16'h001c; // 0x36c8
	13'h1b65: q0 = 16'h6000; // 0x36ca
	13'h1b66: q0 = 16'hfd8e; // 0x36cc
	13'h1b67: q0 = 16'h4a9f; // 0x36ce
	13'h1b68: q0 = 16'h4cdf; // 0x36d0
	13'h1b69: q0 = 16'h20f0; // 0x36d2
	13'h1b6a: q0 = 16'h4e5e; // 0x36d4
	13'h1b6b: q0 = 16'h4e75; // 0x36d6
	13'h1b6c: q0 = 16'h4e56; // 0x36d8
	13'h1b6d: q0 = 16'h0000; // 0x36da
	13'h1b6e: q0 = 16'h48e7; // 0x36dc
	13'h1b6f: q0 = 16'h3f0c; // 0x36de
	13'h1b70: q0 = 16'h2a6e; // 0x36e0
	13'h1b71: q0 = 16'h000c; // 0x36e2
	13'h1b72: q0 = 16'h4245; // 0x36e4
	13'h1b73: q0 = 16'h287c; // 0x36e6
	13'h1b74: q0 = 16'h0001; // 0x36e8
	13'h1b75: q0 = 16'h7bda; // 0x36ea
	13'h1b76: q0 = 16'h4247; // 0x36ec
	13'h1b77: q0 = 16'hbe79; // 0x36ee
	13'h1b78: q0 = 16'h0001; // 0x36f0
	13'h1b79: q0 = 16'h86d6; // 0x36f2
	13'h1b7a: q0 = 16'h6c00; // 0x36f4
	13'h1b7b: q0 = 16'h00b4; // 0x36f6
	13'h1b7c: q0 = 16'h4a6c; // 0x36f8
	13'h1b7d: q0 = 16'h0008; // 0x36fa
	13'h1b7e: q0 = 16'h6702; // 0x36fc
	13'h1b7f: q0 = 16'h5247; // 0x36fe
	13'h1b80: q0 = 16'h0c6c; // 0x3700
	13'h1b81: q0 = 16'h0002; // 0x3702
	13'h1b82: q0 = 16'h0008; // 0x3704
	13'h1b83: q0 = 16'h6600; // 0x3706
	13'h1b84: q0 = 16'h0098; // 0x3708
	13'h1b85: q0 = 16'hbbec; // 0x370a
	13'h1b86: q0 = 16'h000e; // 0x370c
	13'h1b87: q0 = 16'h6700; // 0x370e
	13'h1b88: q0 = 16'h0090; // 0x3710
	13'h1b89: q0 = 16'h302e; // 0x3712
	13'h1b8a: q0 = 16'h0008; // 0x3714
	13'h1b8b: q0 = 16'h226c; // 0x3716
	13'h1b8c: q0 = 16'h0012; // 0x3718
	13'h1b8d: q0 = 16'h9051; // 0x371a
	13'h1b8e: q0 = 16'h3800; // 0x371c
	13'h1b8f: q0 = 16'h4a44; // 0x371e
	13'h1b90: q0 = 16'h6c06; // 0x3720
	13'h1b91: q0 = 16'h3004; // 0x3722
	13'h1b92: q0 = 16'h4440; // 0x3724
	13'h1b93: q0 = 16'h3800; // 0x3726
	13'h1b94: q0 = 16'h302e; // 0x3728
	13'h1b95: q0 = 16'h000a; // 0x372a
	13'h1b96: q0 = 16'h226c; // 0x372c
	13'h1b97: q0 = 16'h0012; // 0x372e
	13'h1b98: q0 = 16'h9069; // 0x3730
	13'h1b99: q0 = 16'h0002; // 0x3732
	13'h1b9a: q0 = 16'h3600; // 0x3734
	13'h1b9b: q0 = 16'h4a43; // 0x3736
	13'h1b9c: q0 = 16'h6c06; // 0x3738
	13'h1b9d: q0 = 16'h3003; // 0x373a
	13'h1b9e: q0 = 16'h4440; // 0x373c
	13'h1b9f: q0 = 16'h3600; // 0x373e
	13'h1ba0: q0 = 16'h200d; // 0x3740
	13'h1ba1: q0 = 16'h6614; // 0x3742
	13'h1ba2: q0 = 16'hb87c; // 0x3744
	13'h1ba3: q0 = 16'h0a00; // 0x3746
	13'h1ba4: q0 = 16'h6c0e; // 0x3748
	13'h1ba5: q0 = 16'hb67c; // 0x374a
	13'h1ba6: q0 = 16'h0a00; // 0x374c
	13'h1ba7: q0 = 16'h6c08; // 0x374e
	13'h1ba8: q0 = 16'h5279; // 0x3750
	13'h1ba9: q0 = 16'h0001; // 0x3752
	13'h1baa: q0 = 16'h7f22; // 0x3754
	13'h1bab: q0 = 16'h7a01; // 0x3756
	13'h1bac: q0 = 16'h4a79; // 0x3758
	13'h1bad: q0 = 16'h0001; // 0x375a
	13'h1bae: q0 = 16'h7f20; // 0x375c
	13'h1baf: q0 = 16'h6706; // 0x375e
	13'h1bb0: q0 = 16'h3c3c; // 0x3760
	13'h1bb1: q0 = 16'h0380; // 0x3762
	13'h1bb2: q0 = 16'h6004; // 0x3764
	13'h1bb3: q0 = 16'h3c2c; // 0x3766
	13'h1bb4: q0 = 16'h0006; // 0x3768
	13'h1bb5: q0 = 16'hb846; // 0x376a
	13'h1bb6: q0 = 16'h6c32; // 0x376c
	13'h1bb7: q0 = 16'hb646; // 0x376e
	13'h1bb8: q0 = 16'h6c2e; // 0x3770
	13'h1bb9: q0 = 16'h206e; // 0x3772
	13'h1bba: q0 = 16'h0010; // 0x3774
	13'h1bbb: q0 = 16'h30ac; // 0x3776
	13'h1bbc: q0 = 16'h000a; // 0x3778
	13'h1bbd: q0 = 16'h206e; // 0x377a
	13'h1bbe: q0 = 16'h0014; // 0x377c
	13'h1bbf: q0 = 16'h30ac; // 0x377e
	13'h1bc0: q0 = 16'h000c; // 0x3780
	13'h1bc1: q0 = 16'h206e; // 0x3782
	13'h1bc2: q0 = 16'h0018; // 0x3784
	13'h1bc3: q0 = 16'h3094; // 0x3786
	13'h1bc4: q0 = 16'h206e; // 0x3788
	13'h1bc5: q0 = 16'h001c; // 0x378a
	13'h1bc6: q0 = 16'h30ac; // 0x378c
	13'h1bc7: q0 = 16'h0002; // 0x378e
	13'h1bc8: q0 = 16'h200d; // 0x3790
	13'h1bc9: q0 = 16'h6708; // 0x3792
	13'h1bca: q0 = 16'h2e8c; // 0x3794
	13'h1bcb: q0 = 16'h4eb9; // 0x3796
	13'h1bcc: q0 = 16'h0000; // 0x3798
	13'h1bcd: q0 = 16'h3a1e; // 0x379a
	13'h1bce: q0 = 16'h200c; // 0x379c
	13'h1bcf: q0 = 16'h603c; // 0x379e
	13'h1bd0: q0 = 16'hd9fc; // 0x37a0
	13'h1bd1: q0 = 16'h0000; // 0x37a2
	13'h1bd2: q0 = 16'h001c; // 0x37a4
	13'h1bd3: q0 = 16'h6000; // 0x37a6
	13'h1bd4: q0 = 16'hff46; // 0x37a8
	13'h1bd5: q0 = 16'h4a45; // 0x37aa
	13'h1bd6: q0 = 16'h6714; // 0x37ac
	13'h1bd7: q0 = 16'h4a79; // 0x37ae
	13'h1bd8: q0 = 16'h0001; // 0x37b0
	13'h1bd9: q0 = 16'h806c; // 0x37b2
	13'h1bda: q0 = 16'h660c; // 0x37b4
	13'h1bdb: q0 = 16'h2ebc; // 0x37b6
	13'h1bdc: q0 = 16'h0000; // 0x37b8
	13'h1bdd: q0 = 16'hc486; // 0x37ba
	13'h1bde: q0 = 16'h4eb9; // 0x37bc
	13'h1bdf: q0 = 16'h0000; // 0x37be
	13'h1be0: q0 = 16'h7dd8; // 0x37c0
	13'h1be1: q0 = 16'h4a45; // 0x37c2
	13'h1be2: q0 = 16'h670a; // 0x37c4
	13'h1be3: q0 = 16'h33fc; // 0x37c6
	13'h1be4: q0 = 16'h0001; // 0x37c8
	13'h1be5: q0 = 16'h0001; // 0x37ca
	13'h1be6: q0 = 16'h806c; // 0x37cc
	13'h1be7: q0 = 16'h600a; // 0x37ce
	13'h1be8: q0 = 16'h200d; // 0x37d0
	13'h1be9: q0 = 16'h6606; // 0x37d2
	13'h1bea: q0 = 16'h4279; // 0x37d4
	13'h1beb: q0 = 16'h0001; // 0x37d6
	13'h1bec: q0 = 16'h806c; // 0x37d8
	13'h1bed: q0 = 16'h7000; // 0x37da
	13'h1bee: q0 = 16'h4a9f; // 0x37dc
	13'h1bef: q0 = 16'h4cdf; // 0x37de
	13'h1bf0: q0 = 16'h30f8; // 0x37e0
	13'h1bf1: q0 = 16'h4e5e; // 0x37e2
	13'h1bf2: q0 = 16'h4e75; // 0x37e4
	13'h1bf3: q0 = 16'h4e56; // 0x37e6
	13'h1bf4: q0 = 16'h0000; // 0x37e8
	13'h1bf5: q0 = 16'h48e7; // 0x37ea
	13'h1bf6: q0 = 16'h3f0c; // 0x37ec
	13'h1bf7: q0 = 16'h3e2e; // 0x37ee
	13'h1bf8: q0 = 16'h0008; // 0x37f0
	13'h1bf9: q0 = 16'h3c2e; // 0x37f2
	13'h1bfa: q0 = 16'h000a; // 0x37f4
	13'h1bfb: q0 = 16'h0c79; // 0x37f6
	13'h1bfc: q0 = 16'h001a; // 0x37f8
	13'h1bfd: q0 = 16'h0001; // 0x37fa
	13'h1bfe: q0 = 16'h86d6; // 0x37fc
	13'h1bff: q0 = 16'h660e; // 0x37fe
	13'h1c00: q0 = 16'h4a79; // 0x3800
	13'h1c01: q0 = 16'h0001; // 0x3802
	13'h1c02: q0 = 16'h7bd6; // 0x3804
	13'h1c03: q0 = 16'h6706; // 0x3806
	13'h1c04: q0 = 16'h7000; // 0x3808
	13'h1c05: q0 = 16'h6000; // 0x380a
	13'h1c06: q0 = 16'h00c2; // 0x380c
	13'h1c07: q0 = 16'h3e86; // 0x380e
	13'h1c08: q0 = 16'h3f07; // 0x3810
	13'h1c09: q0 = 16'h4eb9; // 0x3812
	13'h1c0a: q0 = 16'h0000; // 0x3814
	13'h1c0b: q0 = 16'h82ce; // 0x3816
	13'h1c0c: q0 = 16'h4a5f; // 0x3818
	13'h1c0d: q0 = 16'h3a00; // 0x381a
	13'h1c0e: q0 = 16'h4a45; // 0x381c
	13'h1c0f: q0 = 16'h6606; // 0x381e
	13'h1c10: q0 = 16'h7000; // 0x3820
	13'h1c11: q0 = 16'h6000; // 0x3822
	13'h1c12: q0 = 16'h00aa; // 0x3824
	13'h1c13: q0 = 16'h363c; // 0x3826
	13'h1c14: q0 = 16'h03e7; // 0x3828
	13'h1c15: q0 = 16'h2a7c; // 0x382a
	13'h1c16: q0 = 16'h0001; // 0x382c
	13'h1c17: q0 = 16'h7bda; // 0x382e
	13'h1c18: q0 = 16'h4244; // 0x3830
	13'h1c19: q0 = 16'hb87c; // 0x3832
	13'h1c1a: q0 = 16'h001a; // 0x3834
	13'h1c1b: q0 = 16'h6c26; // 0x3836
	13'h1c1c: q0 = 16'h4a6d; // 0x3838
	13'h1c1d: q0 = 16'h0008; // 0x383a
	13'h1c1e: q0 = 16'h6720; // 0x383c
	13'h1c1f: q0 = 16'h0c6d; // 0x383e
	13'h1c20: q0 = 16'h0002; // 0x3840
	13'h1c21: q0 = 16'h0008; // 0x3842
	13'h1c22: q0 = 16'h660e; // 0x3844
	13'h1c23: q0 = 16'h302d; // 0x3846
	13'h1c24: q0 = 16'h0004; // 0x3848
	13'h1c25: q0 = 16'hb043; // 0x384a
	13'h1c26: q0 = 16'h6c06; // 0x384c
	13'h1c27: q0 = 16'h362d; // 0x384e
	13'h1c28: q0 = 16'h0004; // 0x3850
	13'h1c29: q0 = 16'h284d; // 0x3852
	13'h1c2a: q0 = 16'hdbfc; // 0x3854
	13'h1c2b: q0 = 16'h0000; // 0x3856
	13'h1c2c: q0 = 16'h001c; // 0x3858
	13'h1c2d: q0 = 16'h5244; // 0x385a
	13'h1c2e: q0 = 16'h60d4; // 0x385c
	13'h1c2f: q0 = 16'hb87c; // 0x385e
	13'h1c30: q0 = 16'h001a; // 0x3860
	13'h1c31: q0 = 16'h6604; // 0x3862
	13'h1c32: q0 = 16'h2a4c; // 0x3864
	13'h1c33: q0 = 16'h6006; // 0x3866
	13'h1c34: q0 = 16'h5279; // 0x3868
	13'h1c35: q0 = 16'h0001; // 0x386a
	13'h1c36: q0 = 16'h86d6; // 0x386c
	13'h1c37: q0 = 16'h3005; // 0x386e
	13'h1c38: q0 = 16'h5340; // 0x3870
	13'h1c39: q0 = 16'he740; // 0x3872
	13'h1c3a: q0 = 16'h48c0; // 0x3874
	13'h1c3b: q0 = 16'hd0bc; // 0x3876
	13'h1c3c: q0 = 16'h0000; // 0x3878
	13'h1c3d: q0 = 16'hc9ca; // 0x387a
	13'h1c3e: q0 = 16'h2b40; // 0x387c
	13'h1c3f: q0 = 16'h0016; // 0x387e
	13'h1c40: q0 = 16'h4a6e; // 0x3880
	13'h1c41: q0 = 16'h000c; // 0x3882
	13'h1c42: q0 = 16'h671c; // 0x3884
	13'h1c43: q0 = 16'h206d; // 0x3886
	13'h1c44: q0 = 16'h0012; // 0x3888
	13'h1c45: q0 = 16'h226d; // 0x388a
	13'h1c46: q0 = 16'h0016; // 0x388c
	13'h1c47: q0 = 16'h3151; // 0x388e
	13'h1c48: q0 = 16'h0004; // 0x3890
	13'h1c49: q0 = 16'h206d; // 0x3892
	13'h1c4a: q0 = 16'h0012; // 0x3894
	13'h1c4b: q0 = 16'h226d; // 0x3896
	13'h1c4c: q0 = 16'h0016; // 0x3898
	13'h1c4d: q0 = 16'h3169; // 0x389a
	13'h1c4e: q0 = 16'h0002; // 0x389c
	13'h1c4f: q0 = 16'h0006; // 0x389e
	13'h1c50: q0 = 16'h6012; // 0x38a0
	13'h1c51: q0 = 16'h206d; // 0x38a2
	13'h1c52: q0 = 16'h0012; // 0x38a4
	13'h1c53: q0 = 16'h317c; // 0x38a6
	13'h1c54: q0 = 16'h0030; // 0x38a8
	13'h1c55: q0 = 16'h0004; // 0x38aa
	13'h1c56: q0 = 16'h206d; // 0x38ac
	13'h1c57: q0 = 16'h0012; // 0x38ae
	13'h1c58: q0 = 16'h4268; // 0x38b0
	13'h1c59: q0 = 16'h0006; // 0x38b2
	13'h1c5a: q0 = 16'h206d; // 0x38b4
	13'h1c5b: q0 = 16'h0012; // 0x38b6
	13'h1c5c: q0 = 16'h3087; // 0x38b8
	13'h1c5d: q0 = 16'h206d; // 0x38ba
	13'h1c5e: q0 = 16'h0012; // 0x38bc
	13'h1c5f: q0 = 16'h3146; // 0x38be
	13'h1c60: q0 = 16'h0002; // 0x38c0
	13'h1c61: q0 = 16'h3b7c; // 0x38c2
	13'h1c62: q0 = 16'h0001; // 0x38c4
	13'h1c63: q0 = 16'h0008; // 0x38c6
	13'h1c64: q0 = 16'h3b45; // 0x38c8
	13'h1c65: q0 = 16'h000a; // 0x38ca
	13'h1c66: q0 = 16'h200d; // 0x38cc
	13'h1c67: q0 = 16'h4a9f; // 0x38ce
	13'h1c68: q0 = 16'h4cdf; // 0x38d0
	13'h1c69: q0 = 16'h30f8; // 0x38d2
	13'h1c6a: q0 = 16'h4e5e; // 0x38d4
	13'h1c6b: q0 = 16'h4e75; // 0x38d6
	13'h1c6c: q0 = 16'h4e56; // 0x38d8
	13'h1c6d: q0 = 16'hfffc; // 0x38da
	13'h1c6e: q0 = 16'h48e7; // 0x38dc
	13'h1c6f: q0 = 16'h0f04; // 0x38de
	13'h1c70: q0 = 16'h3e2e; // 0x38e0
	13'h1c71: q0 = 16'h000a; // 0x38e2
	13'h1c72: q0 = 16'h3c2e; // 0x38e4
	13'h1c73: q0 = 16'h000c; // 0x38e6
	13'h1c74: q0 = 16'h42ae; // 0x38e8
	13'h1c75: q0 = 16'hfffc; // 0x38ea
	13'h1c76: q0 = 16'h2a7c; // 0x38ec
	13'h1c77: q0 = 16'h0001; // 0x38ee
	13'h1c78: q0 = 16'h7bda; // 0x38f0
	13'h1c79: q0 = 16'h4245; // 0x38f2
	13'h1c7a: q0 = 16'hba7c; // 0x38f4
	13'h1c7b: q0 = 16'h001a; // 0x38f6
	13'h1c7c: q0 = 16'h6c1c; // 0x38f8
	13'h1c7d: q0 = 16'h4a6d; // 0x38fa
	13'h1c7e: q0 = 16'h0008; // 0x38fc
	13'h1c7f: q0 = 16'h6716; // 0x38fe
	13'h1c80: q0 = 16'h0c6d; // 0x3900
	13'h1c81: q0 = 16'h0005; // 0x3902
	13'h1c82: q0 = 16'h0008; // 0x3904
	13'h1c83: q0 = 16'h6604; // 0x3906
	13'h1c84: q0 = 16'h2d4d; // 0x3908
	13'h1c85: q0 = 16'hfffc; // 0x390a
	13'h1c86: q0 = 16'hdbfc; // 0x390c
	13'h1c87: q0 = 16'h0000; // 0x390e
	13'h1c88: q0 = 16'h001c; // 0x3910
	13'h1c89: q0 = 16'h5245; // 0x3912
	13'h1c8a: q0 = 16'h60de; // 0x3914
	13'h1c8b: q0 = 16'hba7c; // 0x3916
	13'h1c8c: q0 = 16'h001a; // 0x3918
	13'h1c8d: q0 = 16'h6612; // 0x391a
	13'h1c8e: q0 = 16'h4aae; // 0x391c
	13'h1c8f: q0 = 16'hfffc; // 0x391e
	13'h1c90: q0 = 16'h6606; // 0x3920
	13'h1c91: q0 = 16'h7000; // 0x3922
	13'h1c92: q0 = 16'h6058; // 0x3924
	13'h1c93: q0 = 16'h6004; // 0x3926
	13'h1c94: q0 = 16'h2a6e; // 0x3928
	13'h1c95: q0 = 16'hfffc; // 0x392a
	13'h1c96: q0 = 16'h6006; // 0x392c
	13'h1c97: q0 = 16'h5279; // 0x392e
	13'h1c98: q0 = 16'h0001; // 0x3930
	13'h1c99: q0 = 16'h86d6; // 0x3932
	13'h1c9a: q0 = 16'h302e; // 0x3934
	13'h1c9b: q0 = 16'h0008; // 0x3936
	13'h1c9c: q0 = 16'h5340; // 0x3938
	13'h1c9d: q0 = 16'he740; // 0x393a
	13'h1c9e: q0 = 16'h48c0; // 0x393c
	13'h1c9f: q0 = 16'hd0bc; // 0x393e
	13'h1ca0: q0 = 16'h0000; // 0x3940
	13'h1ca1: q0 = 16'hc9ca; // 0x3942
	13'h1ca2: q0 = 16'h2b40; // 0x3944
	13'h1ca3: q0 = 16'h0016; // 0x3946
	13'h1ca4: q0 = 16'h206d; // 0x3948
	13'h1ca5: q0 = 16'h0012; // 0x394a
	13'h1ca6: q0 = 16'h226d; // 0x394c
	13'h1ca7: q0 = 16'h0016; // 0x394e
	13'h1ca8: q0 = 16'h3151; // 0x3950
	13'h1ca9: q0 = 16'h0004; // 0x3952
	13'h1caa: q0 = 16'h206d; // 0x3954
	13'h1cab: q0 = 16'h0012; // 0x3956
	13'h1cac: q0 = 16'h226d; // 0x3958
	13'h1cad: q0 = 16'h0016; // 0x395a
	13'h1cae: q0 = 16'h3169; // 0x395c
	13'h1caf: q0 = 16'h0002; // 0x395e
	13'h1cb0: q0 = 16'h0006; // 0x3960
	13'h1cb1: q0 = 16'h206d; // 0x3962
	13'h1cb2: q0 = 16'h0012; // 0x3964
	13'h1cb3: q0 = 16'h3087; // 0x3966
	13'h1cb4: q0 = 16'h206d; // 0x3968
	13'h1cb5: q0 = 16'h0012; // 0x396a
	13'h1cb6: q0 = 16'h3146; // 0x396c
	13'h1cb7: q0 = 16'h0002; // 0x396e
	13'h1cb8: q0 = 16'h3b7c; // 0x3970
	13'h1cb9: q0 = 16'h0001; // 0x3972
	13'h1cba: q0 = 16'h0008; // 0x3974
	13'h1cbb: q0 = 16'h3b6e; // 0x3976
	13'h1cbc: q0 = 16'h0008; // 0x3978
	13'h1cbd: q0 = 16'h000a; // 0x397a
	13'h1cbe: q0 = 16'h200d; // 0x397c
	13'h1cbf: q0 = 16'h4a9f; // 0x397e
	13'h1cc0: q0 = 16'h4cdf; // 0x3980
	13'h1cc1: q0 = 16'h20e0; // 0x3982
	13'h1cc2: q0 = 16'h4e5e; // 0x3984
	13'h1cc3: q0 = 16'h4e75; // 0x3986
	13'h1cc4: q0 = 16'h4e56; // 0x3988
	13'h1cc5: q0 = 16'h0000; // 0x398a
	13'h1cc6: q0 = 16'h48e7; // 0x398c
	13'h1cc7: q0 = 16'h0104; // 0x398e
	13'h1cc8: q0 = 16'h2a6e; // 0x3990
	13'h1cc9: q0 = 16'h0008; // 0x3992
	13'h1cca: q0 = 16'h3aae; // 0x3994
	13'h1ccb: q0 = 16'h000c; // 0x3996
	13'h1ccc: q0 = 16'h3b6e; // 0x3998
	13'h1ccd: q0 = 16'h000e; // 0x399a
	13'h1cce: q0 = 16'h0002; // 0x399c
	13'h1ccf: q0 = 16'h4a79; // 0x399e
	13'h1cd0: q0 = 16'h0001; // 0x39a0
	13'h1cd1: q0 = 16'h7bd6; // 0x39a2
	13'h1cd2: q0 = 16'h6708; // 0x39a4
	13'h1cd3: q0 = 16'h3b7c; // 0x39a6
	13'h1cd4: q0 = 16'h0700; // 0x39a8
	13'h1cd5: q0 = 16'h0006; // 0x39aa
	13'h1cd6: q0 = 16'h6016; // 0x39ac
	13'h1cd7: q0 = 16'h4a79; // 0x39ae
	13'h1cd8: q0 = 16'h0001; // 0x39b0
	13'h1cd9: q0 = 16'h7f2a; // 0x39b2
	13'h1cda: q0 = 16'h6708; // 0x39b4
	13'h1cdb: q0 = 16'h3b7c; // 0x39b6
	13'h1cdc: q0 = 16'h0400; // 0x39b8
	13'h1cdd: q0 = 16'h0006; // 0x39ba
	13'h1cde: q0 = 16'h6006; // 0x39bc
	13'h1cdf: q0 = 16'h3b7c; // 0x39be
	13'h1ce0: q0 = 16'h0180; // 0x39c0
	13'h1ce1: q0 = 16'h0006; // 0x39c2
	13'h1ce2: q0 = 16'h3b6e; // 0x39c4
	13'h1ce3: q0 = 16'h0010; // 0x39c6
	13'h1ce4: q0 = 16'h001a; // 0x39c8
	13'h1ce5: q0 = 16'h3b6e; // 0x39ca
	13'h1ce6: q0 = 16'h0012; // 0x39cc
	13'h1ce7: q0 = 16'h000c; // 0x39ce
	13'h1ce8: q0 = 16'h3b7c; // 0x39d0
	13'h1ce9: q0 = 16'h0002; // 0x39d2
	13'h1cea: q0 = 16'h0008; // 0x39d4
	13'h1ceb: q0 = 16'h0c6d; // 0x39d6
	13'h1cec: q0 = 16'h0001; // 0x39d8
	13'h1ced: q0 = 16'h000a; // 0x39da
	13'h1cee: q0 = 16'h6606; // 0x39dc
	13'h1cef: q0 = 16'h3b7c; // 0x39de
	13'h1cf0: q0 = 16'h7fff; // 0x39e0
	13'h1cf1: q0 = 16'h0004; // 0x39e2
	13'h1cf2: q0 = 16'h0c6d; // 0x39e4
	13'h1cf3: q0 = 16'h0002; // 0x39e6
	13'h1cf4: q0 = 16'h000a; // 0x39e8
	13'h1cf5: q0 = 16'h6628; // 0x39ea
	13'h1cf6: q0 = 16'h202d; // 0x39ec
	13'h1cf7: q0 = 16'h0012; // 0x39ee
	13'h1cf8: q0 = 16'h5c80; // 0x39f0
	13'h1cf9: q0 = 16'h2e80; // 0x39f2
	13'h1cfa: q0 = 16'h202d; // 0x39f4
	13'h1cfb: q0 = 16'h0012; // 0x39f6
	13'h1cfc: q0 = 16'h5880; // 0x39f8
	13'h1cfd: q0 = 16'h2f00; // 0x39fa
	13'h1cfe: q0 = 16'h3f2d; // 0x39fc
	13'h1cff: q0 = 16'h0002; // 0x39fe
	13'h1d00: q0 = 16'h3f15; // 0x3a00
	13'h1d01: q0 = 16'h4eb9; // 0x3a02
	13'h1d02: q0 = 16'h0000; // 0x3a04
	13'h1d03: q0 = 16'h0a1c; // 0x3a06
	13'h1d04: q0 = 16'h4a9f; // 0x3a08
	13'h1d05: q0 = 16'h3f00; // 0x3a0a
	13'h1d06: q0 = 16'h4eb9; // 0x3a0c
	13'h1d07: q0 = 16'h0000; // 0x3a0e
	13'h1d08: q0 = 16'h3f1e; // 0x3a10
	13'h1d09: q0 = 16'h5c4f; // 0x3a12
	13'h1d0a: q0 = 16'h4a9f; // 0x3a14
	13'h1d0b: q0 = 16'h4cdf; // 0x3a16
	13'h1d0c: q0 = 16'h2000; // 0x3a18
	13'h1d0d: q0 = 16'h4e5e; // 0x3a1a
	13'h1d0e: q0 = 16'h4e75; // 0x3a1c
	13'h1d0f: q0 = 16'h4e56; // 0x3a1e
	13'h1d10: q0 = 16'h0000; // 0x3a20
	13'h1d11: q0 = 16'h48e7; // 0x3a22
	13'h1d12: q0 = 16'h0104; // 0x3a24
	13'h1d13: q0 = 16'h2a6e; // 0x3a26
	13'h1d14: q0 = 16'h0008; // 0x3a28
	13'h1d15: q0 = 16'h3b7c; // 0x3a2a
	13'h1d16: q0 = 16'h0003; // 0x3a2c
	13'h1d17: q0 = 16'h0008; // 0x3a2e
	13'h1d18: q0 = 16'h206d; // 0x3a30
	13'h1d19: q0 = 16'h0012; // 0x3a32
	13'h1d1a: q0 = 16'h322d; // 0x3a34
	13'h1d1b: q0 = 16'h000a; // 0x3a36
	13'h1d1c: q0 = 16'h5341; // 0x3a38
	13'h1d1d: q0 = 16'he341; // 0x3a3a
	13'h1d1e: q0 = 16'h48c1; // 0x3a3c
	13'h1d1f: q0 = 16'hd2bc; // 0x3a3e
	13'h1d20: q0 = 16'h0000; // 0x3a40
	13'h1d21: q0 = 16'hc9c0; // 0x3a42
	13'h1d22: q0 = 16'h2241; // 0x3a44
	13'h1d23: q0 = 16'h3151; // 0x3a46
	13'h1d24: q0 = 16'h0006; // 0x3a48
	13'h1d25: q0 = 16'h0c6d; // 0x3a4a
	13'h1d26: q0 = 16'h0003; // 0x3a4c
	13'h1d27: q0 = 16'h000a; // 0x3a4e
	13'h1d28: q0 = 16'h660e; // 0x3a50
	13'h1d29: q0 = 16'h206d; // 0x3a52
	13'h1d2a: q0 = 16'h0012; // 0x3a54
	13'h1d2b: q0 = 16'h3179; // 0x3a56
	13'h1d2c: q0 = 16'h0000; // 0x3a58
	13'h1d2d: q0 = 16'hc988; // 0x3a5a
	13'h1d2e: q0 = 16'h0004; // 0x3a5c
	13'h1d2f: q0 = 16'h600c; // 0x3a5e
	13'h1d30: q0 = 16'h206d; // 0x3a60
	13'h1d31: q0 = 16'h0012; // 0x3a62
	13'h1d32: q0 = 16'h3179; // 0x3a64
	13'h1d33: q0 = 16'h0000; // 0x3a66
	13'h1d34: q0 = 16'hc99e; // 0x3a68
	13'h1d35: q0 = 16'h0004; // 0x3a6a
	13'h1d36: q0 = 16'h3b7c; // 0x3a6c
	13'h1d37: q0 = 16'h0004; // 0x3a6e
	13'h1d38: q0 = 16'h0004; // 0x3a70
	13'h1d39: q0 = 16'h4a9f; // 0x3a72
	13'h1d3a: q0 = 16'h4cdf; // 0x3a74
	13'h1d3b: q0 = 16'h2000; // 0x3a76
	13'h1d3c: q0 = 16'h4e5e; // 0x3a78
	13'h1d3d: q0 = 16'h4e75; // 0x3a7a
	13'h1d3e: q0 = 16'h4e56; // 0x3a7c
	13'h1d3f: q0 = 16'h0000; // 0x3a7e
	13'h1d40: q0 = 16'h48e7; // 0x3a80
	13'h1d41: q0 = 16'h0f0c; // 0x3a82
	13'h1d42: q0 = 16'h2a6e; // 0x3a84
	13'h1d43: q0 = 16'h0008; // 0x3a86
	13'h1d44: q0 = 16'h287c; // 0x3a88
	13'h1d45: q0 = 16'h0001; // 0x3a8a
	13'h1d46: q0 = 16'h7bda; // 0x3a8c
	13'h1d47: q0 = 16'h4247; // 0x3a8e
	13'h1d48: q0 = 16'hbe7c; // 0x3a90
	13'h1d49: q0 = 16'h001a; // 0x3a92
	13'h1d4a: q0 = 16'h6c00; // 0x3a94
	13'h1d4b: q0 = 16'h0086; // 0x3a96
	13'h1d4c: q0 = 16'hb9cd; // 0x3a98
	13'h1d4d: q0 = 16'h6650; // 0x3a9a
	13'h1d4e: q0 = 16'h4a79; // 0x3a9c
	13'h1d4f: q0 = 16'h0001; // 0x3a9e
	13'h1d50: q0 = 16'h8676; // 0x3aa0
	13'h1d51: q0 = 16'h6724; // 0x3aa2
	13'h1d52: q0 = 16'h397c; // 0x3aa4
	13'h1d53: q0 = 16'h0001; // 0x3aa6
	13'h1d54: q0 = 16'h0008; // 0x3aa8
	13'h1d55: q0 = 16'h3979; // 0x3aaa
	13'h1d56: q0 = 16'h0001; // 0x3aac
	13'h1d57: q0 = 16'h7fa0; // 0x3aae
	13'h1d58: q0 = 16'h000a; // 0x3ab0
	13'h1d59: q0 = 16'h302c; // 0x3ab2
	13'h1d5a: q0 = 16'h000a; // 0x3ab4
	13'h1d5b: q0 = 16'h5340; // 0x3ab6
	13'h1d5c: q0 = 16'he740; // 0x3ab8
	13'h1d5d: q0 = 16'h48c0; // 0x3aba
	13'h1d5e: q0 = 16'hd0bc; // 0x3abc
	13'h1d5f: q0 = 16'h0000; // 0x3abe
	13'h1d60: q0 = 16'hc9ca; // 0x3ac0
	13'h1d61: q0 = 16'h2940; // 0x3ac2
	13'h1d62: q0 = 16'h0016; // 0x3ac4
	13'h1d63: q0 = 16'h6008; // 0x3ac6
	13'h1d64: q0 = 16'h33ec; // 0x3ac8
	13'h1d65: q0 = 16'h000a; // 0x3aca
	13'h1d66: q0 = 16'h0001; // 0x3acc
	13'h1d67: q0 = 16'h7fa0; // 0x3ace
	13'h1d68: q0 = 16'h206c; // 0x3ad0
	13'h1d69: q0 = 16'h0012; // 0x3ad2
	13'h1d6a: q0 = 16'h226c; // 0x3ad4
	13'h1d6b: q0 = 16'h0016; // 0x3ad6
	13'h1d6c: q0 = 16'h3151; // 0x3ad8
	13'h1d6d: q0 = 16'h0004; // 0x3ada
	13'h1d6e: q0 = 16'h206c; // 0x3adc
	13'h1d6f: q0 = 16'h0012; // 0x3ade
	13'h1d70: q0 = 16'h226c; // 0x3ae0
	13'h1d71: q0 = 16'h0016; // 0x3ae2
	13'h1d72: q0 = 16'h3169; // 0x3ae4
	13'h1d73: q0 = 16'h0002; // 0x3ae6
	13'h1d74: q0 = 16'h0006; // 0x3ae8
	13'h1d75: q0 = 16'h6024; // 0x3aea
	13'h1d76: q0 = 16'h206c; // 0x3aec
	13'h1d77: q0 = 16'h0012; // 0x3aee
	13'h1d78: q0 = 16'h4250; // 0x3af0
	13'h1d79: q0 = 16'h206c; // 0x3af2
	13'h1d7a: q0 = 16'h0012; // 0x3af4
	13'h1d7b: q0 = 16'h4268; // 0x3af6
	13'h1d7c: q0 = 16'h0002; // 0x3af8
	13'h1d7d: q0 = 16'h206c; // 0x3afa
	13'h1d7e: q0 = 16'h0012; // 0x3afc
	13'h1d7f: q0 = 16'h317c; // 0x3afe
	13'h1d80: q0 = 16'h0030; // 0x3b00
	13'h1d81: q0 = 16'h0004; // 0x3b02
	13'h1d82: q0 = 16'h206c; // 0x3b04
	13'h1d83: q0 = 16'h0012; // 0x3b06
	13'h1d84: q0 = 16'h4268; // 0x3b08
	13'h1d85: q0 = 16'h0006; // 0x3b0a
	13'h1d86: q0 = 16'h426c; // 0x3b0c
	13'h1d87: q0 = 16'h0008; // 0x3b0e
	13'h1d88: q0 = 16'hd9fc; // 0x3b10
	13'h1d89: q0 = 16'h0000; // 0x3b12
	13'h1d8a: q0 = 16'h001c; // 0x3b14
	13'h1d8b: q0 = 16'h5247; // 0x3b16
	13'h1d8c: q0 = 16'h6000; // 0x3b18
	13'h1d8d: q0 = 16'hff76; // 0x3b1a
	13'h1d8e: q0 = 16'h200d; // 0x3b1c
	13'h1d8f: q0 = 16'h6608; // 0x3b1e
	13'h1d90: q0 = 16'h4279; // 0x3b20
	13'h1d91: q0 = 16'h0001; // 0x3b22
	13'h1d92: q0 = 16'h86d6; // 0x3b24
	13'h1d93: q0 = 16'h6008; // 0x3b26
	13'h1d94: q0 = 16'h33fc; // 0x3b28
	13'h1d95: q0 = 16'h0001; // 0x3b2a
	13'h1d96: q0 = 16'h0001; // 0x3b2c
	13'h1d97: q0 = 16'h86d6; // 0x3b2e
	13'h1d98: q0 = 16'h4279; // 0x3b30
	13'h1d99: q0 = 16'h0001; // 0x3b32
	13'h1d9a: q0 = 16'h7ba0; // 0x3b34
	13'h1d9b: q0 = 16'h2079; // 0x3b36
	13'h1d9c: q0 = 16'h0001; // 0x3b38
	13'h1d9d: q0 = 16'h7fb8; // 0x3b3a
	13'h1d9e: q0 = 16'h3a10; // 0x3b3c
	13'h1d9f: q0 = 16'he545; // 0x3b3e
	13'h1da0: q0 = 16'h3c05; // 0x3b40
	13'h1da1: q0 = 16'he346; // 0x3b42
	13'h1da2: q0 = 16'h2079; // 0x3b44
	13'h1da3: q0 = 16'h0001; // 0x3b46
	13'h1da4: q0 = 16'h7fb8; // 0x3b48
	13'h1da5: q0 = 16'h0c50; // 0x3b4a
	13'h1da6: q0 = 16'h0003; // 0x3b4c
	13'h1da7: q0 = 16'h6e08; // 0x3b4e
	13'h1da8: q0 = 16'h33c5; // 0x3b50
	13'h1da9: q0 = 16'h0001; // 0x3b52
	13'h1daa: q0 = 16'h7fd0; // 0x3b54
	13'h1dab: q0 = 16'h601a; // 0x3b56
	13'h1dac: q0 = 16'h3006; // 0x3b58
	13'h1dad: q0 = 16'h9045; // 0x3b5a
	13'h1dae: q0 = 16'h5440; // 0x3b5c
	13'h1daf: q0 = 16'he440; // 0x3b5e
	13'h1db0: q0 = 16'h3239; // 0x3b60
	13'h1db1: q0 = 16'h0001; // 0x3b62
	13'h1db2: q0 = 16'h757e; // 0x3b64
	13'h1db3: q0 = 16'h5341; // 0x3b66
	13'h1db4: q0 = 16'hc1c1; // 0x3b68
	13'h1db5: q0 = 16'hd045; // 0x3b6a
	13'h1db6: q0 = 16'h33c0; // 0x3b6c
	13'h1db7: q0 = 16'h0001; // 0x3b6e
	13'h1db8: q0 = 16'h7fd0; // 0x3b70
	13'h1db9: q0 = 16'h4a9f; // 0x3b72
	13'h1dba: q0 = 16'h4cdf; // 0x3b74
	13'h1dbb: q0 = 16'h30e0; // 0x3b76
	13'h1dbc: q0 = 16'h4e5e; // 0x3b78
	13'h1dbd: q0 = 16'h4e75; // 0x3b7a
	13'h1dbe: q0 = 16'h4e56; // 0x3b7c
	13'h1dbf: q0 = 16'hfffc; // 0x3b7e
	13'h1dc0: q0 = 16'h206e; // 0x3b80
	13'h1dc1: q0 = 16'h0008; // 0x3b82
	13'h1dc2: q0 = 16'h317c; // 0x3b84
	13'h1dc3: q0 = 16'h0001; // 0x3b86
	13'h1dc4: q0 = 16'h0008; // 0x3b88
	13'h1dc5: q0 = 16'h4e5e; // 0x3b8a
	13'h1dc6: q0 = 16'h4e75; // 0x3b8c
	13'h1dc7: q0 = 16'h4e56; // 0x3b8e
	13'h1dc8: q0 = 16'h0000; // 0x3b90
	13'h1dc9: q0 = 16'h48e7; // 0x3b92
	13'h1dca: q0 = 16'h070c; // 0x3b94
	13'h1dcb: q0 = 16'h2a6e; // 0x3b96
	13'h1dcc: q0 = 16'h0008; // 0x3b98
	13'h1dcd: q0 = 16'h3e2e; // 0x3b9a
	13'h1dce: q0 = 16'h000c; // 0x3b9c
	13'h1dcf: q0 = 16'h286e; // 0x3b9e
	13'h1dd0: q0 = 16'h000e; // 0x3ba0
	13'h1dd1: q0 = 16'h3b7c; // 0x3ba2
	13'h1dd2: q0 = 16'h0400; // 0x3ba4
	13'h1dd3: q0 = 16'h0006; // 0x3ba6
	13'h1dd4: q0 = 16'h3b7c; // 0x3ba8
	13'h1dd5: q0 = 16'h0002; // 0x3baa
	13'h1dd6: q0 = 16'h0008; // 0x3bac
	13'h1dd7: q0 = 16'h2b4c; // 0x3bae
	13'h1dd8: q0 = 16'h000e; // 0x3bb0
	13'h1dd9: q0 = 16'h206d; // 0x3bb2
	13'h1dda: q0 = 16'h0012; // 0x3bb4
	13'h1ddb: q0 = 16'h226d; // 0x3bb6
	13'h1ddc: q0 = 16'h0016; // 0x3bb8
	13'h1ddd: q0 = 16'h3169; // 0x3bba
	13'h1dde: q0 = 16'h0002; // 0x3bbc
	13'h1ddf: q0 = 16'h0006; // 0x3bbe
	13'h1de0: q0 = 16'h0c6d; // 0x3bc0
	13'h1de1: q0 = 16'h0002; // 0x3bc2
	13'h1de2: q0 = 16'h000a; // 0x3bc4
	13'h1de3: q0 = 16'h661c; // 0x3bc6
	13'h1de4: q0 = 16'h202d; // 0x3bc8
	13'h1de5: q0 = 16'h0012; // 0x3bca
	13'h1de6: q0 = 16'h5c80; // 0x3bcc
	13'h1de7: q0 = 16'h2e80; // 0x3bce
	13'h1de8: q0 = 16'h202d; // 0x3bd0
	13'h1de9: q0 = 16'h0012; // 0x3bd2
	13'h1dea: q0 = 16'h5880; // 0x3bd4
	13'h1deb: q0 = 16'h2f00; // 0x3bd6
	13'h1dec: q0 = 16'h3f07; // 0x3bd8
	13'h1ded: q0 = 16'h4eb9; // 0x3bda
	13'h1dee: q0 = 16'h0000; // 0x3bdc
	13'h1def: q0 = 16'h3f1e; // 0x3bde
	13'h1df0: q0 = 16'h5c4f; // 0x3be0
	13'h1df1: q0 = 16'h600c; // 0x3be2
	13'h1df2: q0 = 16'h206d; // 0x3be4
	13'h1df3: q0 = 16'h0012; // 0x3be6
	13'h1df4: q0 = 16'h226d; // 0x3be8
	13'h1df5: q0 = 16'h0016; // 0x3bea
	13'h1df6: q0 = 16'h3151; // 0x3bec
	13'h1df7: q0 = 16'h0004; // 0x3bee
	13'h1df8: q0 = 16'h2039; // 0x3bf0
	13'h1df9: q0 = 16'h0000; // 0x3bf2
	13'h1dfa: q0 = 16'hc8d6; // 0x3bf4
	13'h1dfb: q0 = 16'he380; // 0x3bf6
	13'h1dfc: q0 = 16'hb08c; // 0x3bf8
	13'h1dfd: q0 = 16'h660c; // 0x3bfa
	13'h1dfe: q0 = 16'h2079; // 0x3bfc
	13'h1dff: q0 = 16'h0001; // 0x3bfe
	13'h1e00: q0 = 16'h7fb8; // 0x3c00
	13'h1e01: q0 = 16'h3c10; // 0x3c02
	13'h1e02: q0 = 16'he746; // 0x3c04
	13'h1e03: q0 = 16'h6006; // 0x3c06
	13'h1e04: q0 = 16'h3c39; // 0x3c08
	13'h1e05: q0 = 16'h0001; // 0x3c0a
	13'h1e06: q0 = 16'h7fd0; // 0x3c0c
	13'h1e07: q0 = 16'h0c6d; // 0x3c0e
	13'h1e08: q0 = 16'h0005; // 0x3c10
	13'h1e09: q0 = 16'h000a; // 0x3c12
	13'h1e0a: q0 = 16'h6716; // 0x3c14
	13'h1e0b: q0 = 16'h206d; // 0x3c16
	13'h1e0c: q0 = 16'h0016; // 0x3c18
	13'h1e0d: q0 = 16'h3b68; // 0x3c1a
	13'h1e0e: q0 = 16'h0006; // 0x3c1c
	13'h1e0f: q0 = 16'h0004; // 0x3c1e
	13'h1e10: q0 = 16'h206d; // 0x3c20
	13'h1e11: q0 = 16'h0016; // 0x3c22
	13'h1e12: q0 = 16'h3028; // 0x3c24
	13'h1e13: q0 = 16'h0004; // 0x3c26
	13'h1e14: q0 = 16'hdc40; // 0x3c28
	13'h1e15: q0 = 16'h603a; // 0x3c2a
	13'h1e16: q0 = 16'h4a79; // 0x3c2c
	13'h1e17: q0 = 16'h0001; // 0x3c2e
	13'h1e18: q0 = 16'h7f20; // 0x3c30
	13'h1e19: q0 = 16'h670c; // 0x3c32
	13'h1e1a: q0 = 16'h3b7c; // 0x3c34
	13'h1e1b: q0 = 16'h0014; // 0x3c36
	13'h1e1c: q0 = 16'h0004; // 0x3c38
	13'h1e1d: q0 = 16'h3c3c; // 0x3c3a
	13'h1e1e: q0 = 16'h0280; // 0x3c3c
	13'h1e1f: q0 = 16'h6026; // 0x3c3e
	13'h1e20: q0 = 16'h3ebc; // 0x3c40
	13'h1e21: q0 = 16'h00ff; // 0x3c42
	13'h1e22: q0 = 16'h3f3c; // 0x3c44
	13'h1e23: q0 = 16'h0010; // 0x3c46
	13'h1e24: q0 = 16'h4eb9; // 0x3c48
	13'h1e25: q0 = 16'h0000; // 0x3c4a
	13'h1e26: q0 = 16'h8e6c; // 0x3c4c
	13'h1e27: q0 = 16'h4a5f; // 0x3c4e
	13'h1e28: q0 = 16'h3b40; // 0x3c50
	13'h1e29: q0 = 16'h0004; // 0x3c52
	13'h1e2a: q0 = 16'h3ebc; // 0x3c54
	13'h1e2b: q0 = 16'h0280; // 0x3c56
	13'h1e2c: q0 = 16'h3f3c; // 0x3c58
	13'h1e2d: q0 = 16'h0100; // 0x3c5a
	13'h1e2e: q0 = 16'h4eb9; // 0x3c5c
	13'h1e2f: q0 = 16'h0000; // 0x3c5e
	13'h1e30: q0 = 16'h8e6c; // 0x3c60
	13'h1e31: q0 = 16'h4a5f; // 0x3c62
	13'h1e32: q0 = 16'hdc40; // 0x3c64
	13'h1e33: q0 = 16'h3e86; // 0x3c66
	13'h1e34: q0 = 16'h3f07; // 0x3c68
	13'h1e35: q0 = 16'h4eb9; // 0x3c6a
	13'h1e36: q0 = 16'h0000; // 0x3c6c
	13'h1e37: q0 = 16'h1280; // 0x3c6e
	13'h1e38: q0 = 16'h4a5f; // 0x3c70
	13'h1e39: q0 = 16'h3a80; // 0x3c72
	13'h1e3a: q0 = 16'h3e86; // 0x3c74
	13'h1e3b: q0 = 16'h3f07; // 0x3c76
	13'h1e3c: q0 = 16'h4eb9; // 0x3c78
	13'h1e3d: q0 = 16'h0000; // 0x3c7a
	13'h1e3e: q0 = 16'ha730; // 0x3c7c
	13'h1e3f: q0 = 16'h4a5f; // 0x3c7e
	13'h1e40: q0 = 16'h3b40; // 0x3c80
	13'h1e41: q0 = 16'h0002; // 0x3c82
	13'h1e42: q0 = 16'h3b47; // 0x3c84
	13'h1e43: q0 = 16'h000c; // 0x3c86
	13'h1e44: q0 = 16'h4a9f; // 0x3c88
	13'h1e45: q0 = 16'h4cdf; // 0x3c8a
	13'h1e46: q0 = 16'h30c0; // 0x3c8c
	13'h1e47: q0 = 16'h4e5e; // 0x3c8e
	13'h1e48: q0 = 16'h4e75; // 0x3c90
	13'h1e49: q0 = 16'h4e56; // 0x3c92
	13'h1e4a: q0 = 16'h0000; // 0x3c94
	13'h1e4b: q0 = 16'h48e7; // 0x3c96
	13'h1e4c: q0 = 16'h0104; // 0x3c98
	13'h1e4d: q0 = 16'h2a6e; // 0x3c9a
	13'h1e4e: q0 = 16'h0008; // 0x3c9c
	13'h1e4f: q0 = 16'h206d; // 0x3c9e
	13'h1e50: q0 = 16'h0012; // 0x3ca0
	13'h1e51: q0 = 16'h30ae; // 0x3ca2
	13'h1e52: q0 = 16'h000c; // 0x3ca4
	13'h1e53: q0 = 16'h206d; // 0x3ca6
	13'h1e54: q0 = 16'h0012; // 0x3ca8
	13'h1e55: q0 = 16'h316e; // 0x3caa
	13'h1e56: q0 = 16'h000e; // 0x3cac
	13'h1e57: q0 = 16'h0002; // 0x3cae
	13'h1e58: q0 = 16'h4a6e; // 0x3cb0
	13'h1e59: q0 = 16'h0010; // 0x3cb2
	13'h1e5a: q0 = 16'h671a; // 0x3cb4
	13'h1e5b: q0 = 16'h206d; // 0x3cb6
	13'h1e5c: q0 = 16'h0012; // 0x3cb8
	13'h1e5d: q0 = 16'h226d; // 0x3cba
	13'h1e5e: q0 = 16'h0016; // 0x3cbc
	13'h1e5f: q0 = 16'h3151; // 0x3cbe
	13'h1e60: q0 = 16'h0004; // 0x3cc0
	13'h1e61: q0 = 16'h206d; // 0x3cc2
	13'h1e62: q0 = 16'h0012; // 0x3cc4
	13'h1e63: q0 = 16'h226d; // 0x3cc6
	13'h1e64: q0 = 16'h0016; // 0x3cc8
	13'h1e65: q0 = 16'h3169; // 0x3cca
	13'h1e66: q0 = 16'h0002; // 0x3ccc
	13'h1e67: q0 = 16'h0006; // 0x3cce
	13'h1e68: q0 = 16'h4a9f; // 0x3cd0
	13'h1e69: q0 = 16'h4cdf; // 0x3cd2
	13'h1e6a: q0 = 16'h2000; // 0x3cd4
	13'h1e6b: q0 = 16'h4e5e; // 0x3cd6
	13'h1e6c: q0 = 16'h4e75; // 0x3cd8
	13'h1e6d: q0 = 16'h4e56; // 0x3cda
	13'h1e6e: q0 = 16'h0000; // 0x3cdc
	13'h1e6f: q0 = 16'h48e7; // 0x3cde
	13'h1e70: q0 = 16'h0300; // 0x3ce0
	13'h1e71: q0 = 16'h4247; // 0x3ce2
	13'h1e72: q0 = 16'hbe7c; // 0x3ce4
	13'h1e73: q0 = 16'h000a; // 0x3ce6
	13'h1e74: q0 = 16'h6c24; // 0x3ce8
	13'h1e75: q0 = 16'h3007; // 0x3cea
	13'h1e76: q0 = 16'he340; // 0x3cec
	13'h1e77: q0 = 16'h48c0; // 0x3cee
	13'h1e78: q0 = 16'hd0bc; // 0x3cf0
	13'h1e79: q0 = 16'h0001; // 0x3cf2
	13'h1e7a: q0 = 16'h86b8; // 0x3cf4
	13'h1e7b: q0 = 16'h2040; // 0x3cf6
	13'h1e7c: q0 = 16'h3207; // 0x3cf8
	13'h1e7d: q0 = 16'h48c1; // 0x3cfa
	13'h1e7e: q0 = 16'hd2bc; // 0x3cfc
	13'h1e7f: q0 = 16'h0000; // 0x3cfe
	13'h1e80: q0 = 16'hc8da; // 0x3d00
	13'h1e81: q0 = 16'h2241; // 0x3d02
	13'h1e82: q0 = 16'h1211; // 0x3d04
	13'h1e83: q0 = 16'h4881; // 0x3d06
	13'h1e84: q0 = 16'h3081; // 0x3d08
	13'h1e85: q0 = 16'h5247; // 0x3d0a
	13'h1e86: q0 = 16'h60d6; // 0x3d0c
	13'h1e87: q0 = 16'h4a9f; // 0x3d0e
	13'h1e88: q0 = 16'h4cdf; // 0x3d10
	13'h1e89: q0 = 16'h0080; // 0x3d12
	13'h1e8a: q0 = 16'h4e5e; // 0x3d14
	13'h1e8b: q0 = 16'h4e75; // 0x3d16
	13'h1e8c: q0 = 16'h4e56; // 0x3d18
	13'h1e8d: q0 = 16'h0000; // 0x3d1a
	13'h1e8e: q0 = 16'h48e7; // 0x3d1c
	13'h1e8f: q0 = 16'h1f04; // 0x3d1e
	13'h1e90: q0 = 16'h3e2e; // 0x3d20
	13'h1e91: q0 = 16'h000c; // 0x3d22
	13'h1e92: q0 = 16'h3c2e; // 0x3d24
	13'h1e93: q0 = 16'h000e; // 0x3d26
	13'h1e94: q0 = 16'h3a2e; // 0x3d28
	13'h1e95: q0 = 16'h0008; // 0x3d2a
	13'h1e96: q0 = 16'hca7c; // 0x3d2c
	13'h1e97: q0 = 16'h001f; // 0x3d2e
	13'h1e98: q0 = 16'h4a79; // 0x3d30
	13'h1e99: q0 = 16'h0001; // 0x3d32
	13'h1e9a: q0 = 16'h7fa6; // 0x3d34
	13'h1e9b: q0 = 16'h6706; // 0x3d36
	13'h1e9c: q0 = 16'h701f; // 0x3d38
	13'h1e9d: q0 = 16'h9045; // 0x3d3a
	13'h1e9e: q0 = 16'h3a00; // 0x3d3c
	13'h1e9f: q0 = 16'h4a45; // 0x3d3e
	13'h1ea0: q0 = 16'h6606; // 0x3d40
	13'h1ea1: q0 = 16'h383c; // 0x3d42
	13'h1ea2: q0 = 16'h07c0; // 0x3d44
	13'h1ea3: q0 = 16'h6006; // 0x3d46
	13'h1ea4: q0 = 16'h3805; // 0x3d48
	13'h1ea5: q0 = 16'h5344; // 0x3d4a
	13'h1ea6: q0 = 16'hed44; // 0x3d4c
	13'h1ea7: q0 = 16'h3a2e; // 0x3d4e
	13'h1ea8: q0 = 16'h000a; // 0x3d50
	13'h1ea9: q0 = 16'hca7c; // 0x3d52
	13'h1eaa: q0 = 16'h001f; // 0x3d54
	13'h1eab: q0 = 16'hba7c; // 0x3d56
	13'h1eac: q0 = 16'h0004; // 0x3d58
	13'h1ead: q0 = 16'h6c02; // 0x3d5a
	13'h1eae: q0 = 16'h7a04; // 0x3d5c
	13'h1eaf: q0 = 16'h4a79; // 0x3d5e
	13'h1eb0: q0 = 16'h0001; // 0x3d60
	13'h1eb1: q0 = 16'h7fa6; // 0x3d62
	13'h1eb2: q0 = 16'h6706; // 0x3d64
	13'h1eb3: q0 = 16'h7023; // 0x3d66
	13'h1eb4: q0 = 16'h9045; // 0x3d68
	13'h1eb5: q0 = 16'h3a00; // 0x3d6a
	13'h1eb6: q0 = 16'h701f; // 0x3d6c
	13'h1eb7: q0 = 16'h9045; // 0x3d6e
	13'h1eb8: q0 = 16'he340; // 0x3d70
	13'h1eb9: q0 = 16'hd840; // 0x3d72
	13'h1eba: q0 = 16'h3044; // 0x3d74
	13'h1ebb: q0 = 16'h2a48; // 0x3d76
	13'h1ebc: q0 = 16'hdbf9; // 0x3d78
	13'h1ebd: q0 = 16'h0000; // 0x3d7a
	13'h1ebe: q0 = 16'hc980; // 0x3d7c
	13'h1ebf: q0 = 16'h3006; // 0x3d7e
	13'h1ec0: q0 = 16'hc07c; // 0x3d80
	13'h1ec1: q0 = 16'h003f; // 0x3d82
	13'h1ec2: q0 = 16'he140; // 0x3d84
	13'h1ec3: q0 = 16'h3207; // 0x3d86
	13'h1ec4: q0 = 16'hc27c; // 0x3d88
	13'h1ec5: q0 = 16'h0100; // 0x3d8a
	13'h1ec6: q0 = 16'hef41; // 0x3d8c
	13'h1ec7: q0 = 16'h8041; // 0x3d8e
	13'h1ec8: q0 = 16'h3207; // 0x3d90
	13'h1ec9: q0 = 16'hc27c; // 0x3d92
	13'h1eca: q0 = 16'h00ff; // 0x3d94
	13'h1ecb: q0 = 16'h8041; // 0x3d96
	13'h1ecc: q0 = 16'h3a80; // 0x3d98
	13'h1ecd: q0 = 16'h4a9f; // 0x3d9a
	13'h1ece: q0 = 16'h4cdf; // 0x3d9c
	13'h1ecf: q0 = 16'h20f0; // 0x3d9e
	13'h1ed0: q0 = 16'h4e5e; // 0x3da0
	13'h1ed1: q0 = 16'h4e75; // 0x3da2
	13'h1ed2: q0 = 16'h4e56; // 0x3da4
	13'h1ed3: q0 = 16'hfffc; // 0x3da6
	13'h1ed4: q0 = 16'h23ee; // 0x3da8
	13'h1ed5: q0 = 16'h0008; // 0x3daa
	13'h1ed6: q0 = 16'h0001; // 0x3dac
	13'h1ed7: q0 = 16'h7f60; // 0x3dae
	13'h1ed8: q0 = 16'h4ab9; // 0x3db0
	13'h1ed9: q0 = 16'h0001; // 0x3db2
	13'h1eda: q0 = 16'h7f60; // 0x3db4
	13'h1edb: q0 = 16'h6702; // 0x3db6
	13'h1edc: q0 = 16'h60f6; // 0x3db8
	13'h1edd: q0 = 16'h4e5e; // 0x3dba
	13'h1ede: q0 = 16'h4e75; // 0x3dbc
	13'h1edf: q0 = 16'h4e56; // 0x3dbe
	13'h1ee0: q0 = 16'h0000; // 0x3dc0
	13'h1ee1: q0 = 16'h48e7; // 0x3dc2
	13'h1ee2: q0 = 16'h071c; // 0x3dc4
	13'h1ee3: q0 = 16'h2a6e; // 0x3dc6
	13'h1ee4: q0 = 16'h000c; // 0x3dc8
	13'h1ee5: q0 = 16'h286e; // 0x3dca
	13'h1ee6: q0 = 16'h0010; // 0x3dcc
	13'h1ee7: q0 = 16'h3e2e; // 0x3dce
	13'h1ee8: q0 = 16'h0008; // 0x3dd0
	13'h1ee9: q0 = 16'hee47; // 0x3dd2
	13'h1eea: q0 = 16'he647; // 0x3dd4
	13'h1eeb: q0 = 16'hce7c; // 0x3dd6
	13'h1eec: q0 = 16'h001f; // 0x3dd8
	13'h1eed: q0 = 16'h4a79; // 0x3dda
	13'h1eee: q0 = 16'h0001; // 0x3ddc
	13'h1eef: q0 = 16'h7fa6; // 0x3dde
	13'h1ef0: q0 = 16'h6706; // 0x3de0
	13'h1ef1: q0 = 16'h701f; // 0x3de2
	13'h1ef2: q0 = 16'h9047; // 0x3de4
	13'h1ef3: q0 = 16'h3e00; // 0x3de6
	13'h1ef4: q0 = 16'h4a47; // 0x3de8
	13'h1ef5: q0 = 16'h6606; // 0x3dea
	13'h1ef6: q0 = 16'h3c3c; // 0x3dec
	13'h1ef7: q0 = 16'h07c0; // 0x3dee
	13'h1ef8: q0 = 16'h6006; // 0x3df0
	13'h1ef9: q0 = 16'h3c07; // 0x3df2
	13'h1efa: q0 = 16'h5346; // 0x3df4
	13'h1efb: q0 = 16'hed46; // 0x3df6
	13'h1efc: q0 = 16'h3e2e; // 0x3df8
	13'h1efd: q0 = 16'h000a; // 0x3dfa
	13'h1efe: q0 = 16'hee47; // 0x3dfc
	13'h1eff: q0 = 16'he647; // 0x3dfe
	13'h1f00: q0 = 16'hce7c; // 0x3e00
	13'h1f01: q0 = 16'h001f; // 0x3e02
	13'h1f02: q0 = 16'hbe7c; // 0x3e04
	13'h1f03: q0 = 16'h0004; // 0x3e06
	13'h1f04: q0 = 16'h6c02; // 0x3e08
	13'h1f05: q0 = 16'h7e04; // 0x3e0a
	13'h1f06: q0 = 16'h4a79; // 0x3e0c
	13'h1f07: q0 = 16'h0001; // 0x3e0e
	13'h1f08: q0 = 16'h7fa6; // 0x3e10
	13'h1f09: q0 = 16'h6706; // 0x3e12
	13'h1f0a: q0 = 16'h7023; // 0x3e14
	13'h1f0b: q0 = 16'h9047; // 0x3e16
	13'h1f0c: q0 = 16'h3e00; // 0x3e18
	13'h1f0d: q0 = 16'h701f; // 0x3e1a
	13'h1f0e: q0 = 16'h9047; // 0x3e1c
	13'h1f0f: q0 = 16'he340; // 0x3e1e
	13'h1f10: q0 = 16'hdc40; // 0x3e20
	13'h1f11: q0 = 16'h3046; // 0x3e22
	13'h1f12: q0 = 16'h2648; // 0x3e24
	13'h1f13: q0 = 16'hd7f9; // 0x3e26
	13'h1f14: q0 = 16'h0000; // 0x3e28
	13'h1f15: q0 = 16'hc984; // 0x3e2a
	13'h1f16: q0 = 16'h3013; // 0x3e2c
	13'h1f17: q0 = 16'he040; // 0x3e2e
	13'h1f18: q0 = 16'hc07c; // 0x3e30
	13'h1f19: q0 = 16'h003f; // 0x3e32
	13'h1f1a: q0 = 16'h3880; // 0x3e34
	13'h1f1b: q0 = 16'h3013; // 0x3e36
	13'h1f1c: q0 = 16'hee40; // 0x3e38
	13'h1f1d: q0 = 16'hc07c; // 0x3e3a
	13'h1f1e: q0 = 16'h0100; // 0x3e3c
	13'h1f1f: q0 = 16'h3213; // 0x3e3e
	13'h1f20: q0 = 16'hc27c; // 0x3e40
	13'h1f21: q0 = 16'h00ff; // 0x3e42
	13'h1f22: q0 = 16'h8041; // 0x3e44
	13'h1f23: q0 = 16'h3a80; // 0x3e46
	13'h1f24: q0 = 16'h4a9f; // 0x3e48
	13'h1f25: q0 = 16'h4cdf; // 0x3e4a
	13'h1f26: q0 = 16'h38c0; // 0x3e4c
	13'h1f27: q0 = 16'h4e5e; // 0x3e4e
	13'h1f28: q0 = 16'h4e75; // 0x3e50
	13'h1f29: q0 = 16'h4e56; // 0x3e52
	13'h1f2a: q0 = 16'h0000; // 0x3e54
	13'h1f2b: q0 = 16'h48e7; // 0x3e56
	13'h1f2c: q0 = 16'h0700; // 0x3e58
	13'h1f2d: q0 = 16'h3e2e; // 0x3e5a
	13'h1f2e: q0 = 16'h0008; // 0x3e5c
	13'h1f2f: q0 = 16'h2079; // 0x3e5e
	13'h1f30: q0 = 16'h0001; // 0x3e60
	13'h1f31: q0 = 16'h7fb8; // 0x3e62
	13'h1f32: q0 = 16'h0c50; // 0x3e64
	13'h1f33: q0 = 16'h0005; // 0x3e66
	13'h1f34: q0 = 16'h6c14; // 0x3e68
	13'h1f35: q0 = 16'h3ebc; // 0x3e6a
	13'h1f36: q0 = 16'h0004; // 0x3e6c
	13'h1f37: q0 = 16'h3f3c; // 0x3e6e
	13'h1f38: q0 = 16'h0001; // 0x3e70
	13'h1f39: q0 = 16'h4eb9; // 0x3e72
	13'h1f3a: q0 = 16'h0000; // 0x3e74
	13'h1f3b: q0 = 16'h8e6c; // 0x3e76
	13'h1f3c: q0 = 16'h4a5f; // 0x3e78
	13'h1f3d: q0 = 16'h3c00; // 0x3e7a
	13'h1f3e: q0 = 16'h605c; // 0x3e7c
	13'h1f3f: q0 = 16'hbe7c; // 0x3e7e
	13'h1f40: q0 = 16'h0005; // 0x3e80
	13'h1f41: q0 = 16'h6604; // 0x3e82
	13'h1f42: q0 = 16'h7c05; // 0x3e84
	13'h1f43: q0 = 16'h6052; // 0x3e86
	13'h1f44: q0 = 16'hbe7c; // 0x3e88
	13'h1f45: q0 = 16'h0006; // 0x3e8a
	13'h1f46: q0 = 16'h6604; // 0x3e8c
	13'h1f47: q0 = 16'h7c01; // 0x3e8e
	13'h1f48: q0 = 16'h6048; // 0x3e90
	13'h1f49: q0 = 16'hbe7c; // 0x3e92
	13'h1f4a: q0 = 16'h0008; // 0x3e94
	13'h1f4b: q0 = 16'h6604; // 0x3e96
	13'h1f4c: q0 = 16'h7c03; // 0x3e98
	13'h1f4d: q0 = 16'h603e; // 0x3e9a
	13'h1f4e: q0 = 16'hbe7c; // 0x3e9c
	13'h1f4f: q0 = 16'h0001; // 0x3e9e
	13'h1f50: q0 = 16'h6604; // 0x3ea0
	13'h1f51: q0 = 16'h7c04; // 0x3ea2
	13'h1f52: q0 = 16'h6034; // 0x3ea4
	13'h1f53: q0 = 16'hbe7c; // 0x3ea6
	13'h1f54: q0 = 16'h0003; // 0x3ea8
	13'h1f55: q0 = 16'h6604; // 0x3eaa
	13'h1f56: q0 = 16'h7c02; // 0x3eac
	13'h1f57: q0 = 16'h602a; // 0x3eae
	13'h1f58: q0 = 16'h4a47; // 0x3eb0
	13'h1f59: q0 = 16'h6614; // 0x3eb2
	13'h1f5a: q0 = 16'h3ebc; // 0x3eb4
	13'h1f5b: q0 = 16'h0005; // 0x3eb6
	13'h1f5c: q0 = 16'h3f3c; // 0x3eb8
	13'h1f5d: q0 = 16'h0001; // 0x3eba
	13'h1f5e: q0 = 16'h4eb9; // 0x3ebc
	13'h1f5f: q0 = 16'h0000; // 0x3ebe
	13'h1f60: q0 = 16'h8e6c; // 0x3ec0
	13'h1f61: q0 = 16'h4a5f; // 0x3ec2
	13'h1f62: q0 = 16'h3c00; // 0x3ec4
	13'h1f63: q0 = 16'h6012; // 0x3ec6
	13'h1f64: q0 = 16'h3ebc; // 0x3ec8
	13'h1f65: q0 = 16'h0004; // 0x3eca
	13'h1f66: q0 = 16'h3f3c; // 0x3ecc
	13'h1f67: q0 = 16'h0001; // 0x3ece
	13'h1f68: q0 = 16'h4eb9; // 0x3ed0
	13'h1f69: q0 = 16'h0000; // 0x3ed2
	13'h1f6a: q0 = 16'h8e6c; // 0x3ed4
	13'h1f6b: q0 = 16'h4a5f; // 0x3ed6
	13'h1f6c: q0 = 16'h3c00; // 0x3ed8
	13'h1f6d: q0 = 16'h3006; // 0x3eda
	13'h1f6e: q0 = 16'h4a9f; // 0x3edc
	13'h1f6f: q0 = 16'h4cdf; // 0x3ede
	13'h1f70: q0 = 16'h00c0; // 0x3ee0
	13'h1f71: q0 = 16'h4e5e; // 0x3ee2
	13'h1f72: q0 = 16'h4e75; // 0x3ee4
	13'h1f73: q0 = 16'h4e56; // 0x3ee6
	13'h1f74: q0 = 16'h0000; // 0x3ee8
	13'h1f75: q0 = 16'h48e7; // 0x3eea
	13'h1f76: q0 = 16'h0304; // 0x3eec
	13'h1f77: q0 = 16'h2a6e; // 0x3eee
	13'h1f78: q0 = 16'h0008; // 0x3ef0
	13'h1f79: q0 = 16'h3e2e; // 0x3ef2
	13'h1f7a: q0 = 16'h000c; // 0x3ef4
	13'h1f7b: q0 = 16'hbe7c; // 0x3ef6
	13'h1f7c: q0 = 16'h0012; // 0x3ef8
	13'h1f7d: q0 = 16'h6f10; // 0x3efa
	13'h1f7e: q0 = 16'hbe7c; // 0x3efc
	13'h1f7f: q0 = 16'h0036; // 0x3efe
	13'h1f80: q0 = 16'h6e0a; // 0x3f00
	13'h1f81: q0 = 16'h3015; // 0x3f02
	13'h1f82: q0 = 16'h807c; // 0x3f04
	13'h1f83: q0 = 16'h0080; // 0x3f06
	13'h1f84: q0 = 16'h3a80; // 0x3f08
	13'h1f85: q0 = 16'h6008; // 0x3f0a
	13'h1f86: q0 = 16'h3015; // 0x3f0c
	13'h1f87: q0 = 16'hc07c; // 0x3f0e
	13'h1f88: q0 = 16'h003f; // 0x3f10
	13'h1f89: q0 = 16'h3a80; // 0x3f12
	13'h1f8a: q0 = 16'h4a9f; // 0x3f14
	13'h1f8b: q0 = 16'h4cdf; // 0x3f16
	13'h1f8c: q0 = 16'h2080; // 0x3f18
	13'h1f8d: q0 = 16'h4e5e; // 0x3f1a
	13'h1f8e: q0 = 16'h4e75; // 0x3f1c
	13'h1f8f: q0 = 16'h4e56; // 0x3f1e
	13'h1f90: q0 = 16'h0000; // 0x3f20
	13'h1f91: q0 = 16'h48e7; // 0x3f22
	13'h1f92: q0 = 16'h0300; // 0x3f24
	13'h1f93: q0 = 16'h4247; // 0x3f26
	13'h1f94: q0 = 16'h3007; // 0x3f28
	13'h1f95: q0 = 16'h48c0; // 0x3f2a
	13'h1f96: q0 = 16'hd0bc; // 0x3f2c
	13'h1f97: q0 = 16'h0000; // 0x3f2e
	13'h1f98: q0 = 16'hc9f2; // 0x3f30
	13'h1f99: q0 = 16'h2040; // 0x3f32
	13'h1f9a: q0 = 16'h1010; // 0x3f34
	13'h1f9b: q0 = 16'h4880; // 0x3f36
	13'h1f9c: q0 = 16'hb06e; // 0x3f38
	13'h1f9d: q0 = 16'h0008; // 0x3f3a
	13'h1f9e: q0 = 16'h6e04; // 0x3f3c
	13'h1f9f: q0 = 16'h5247; // 0x3f3e
	13'h1fa0: q0 = 16'h60e6; // 0x3f40
	13'h1fa1: q0 = 16'hbe7c; // 0x3f42
	13'h1fa2: q0 = 16'h0008; // 0x3f44
	13'h1fa3: q0 = 16'h6602; // 0x3f46
	13'h1fa4: q0 = 16'h4247; // 0x3f48
	13'h1fa5: q0 = 16'h206e; // 0x3f4a
	13'h1fa6: q0 = 16'h000a; // 0x3f4c
	13'h1fa7: q0 = 16'h3207; // 0x3f4e
	13'h1fa8: q0 = 16'h48c1; // 0x3f50
	13'h1fa9: q0 = 16'hd2bc; // 0x3f52
	13'h1faa: q0 = 16'h0000; // 0x3f54
	13'h1fab: q0 = 16'hc9fc; // 0x3f56
	13'h1fac: q0 = 16'h2241; // 0x3f58
	13'h1fad: q0 = 16'h1211; // 0x3f5a
	13'h1fae: q0 = 16'h4881; // 0x3f5c
	13'h1faf: q0 = 16'h3081; // 0x3f5e
	13'h1fb0: q0 = 16'h3007; // 0x3f60
	13'h1fb1: q0 = 16'h48c0; // 0x3f62
	13'h1fb2: q0 = 16'hd0bc; // 0x3f64
	13'h1fb3: q0 = 16'h0000; // 0x3f66
	13'h1fb4: q0 = 16'hca04; // 0x3f68
	13'h1fb5: q0 = 16'h2040; // 0x3f6a
	13'h1fb6: q0 = 16'h1010; // 0x3f6c
	13'h1fb7: q0 = 16'h4880; // 0x3f6e
	13'h1fb8: q0 = 16'h226e; // 0x3f70
	13'h1fb9: q0 = 16'h000e; // 0x3f72
	13'h1fba: q0 = 16'h8151; // 0x3f74
	13'h1fbb: q0 = 16'h4a9f; // 0x3f76
	13'h1fbc: q0 = 16'h4cdf; // 0x3f78
	13'h1fbd: q0 = 16'h0080; // 0x3f7a
	13'h1fbe: q0 = 16'h4e5e; // 0x3f7c
	13'h1fbf: q0 = 16'h4e75; // 0x3f7e
	13'h1fc0: q0 = 16'h4e56; // 0x3f80
	13'h1fc1: q0 = 16'hfffc; // 0x3f82
	13'h1fc2: q0 = 16'h3eae; // 0x3f84
	13'h1fc3: q0 = 16'h000e; // 0x3f86
	13'h1fc4: q0 = 16'h3f2e; // 0x3f88
	13'h1fc5: q0 = 16'h000c; // 0x3f8a
	13'h1fc6: q0 = 16'h302e; // 0x3f8c
	13'h1fc7: q0 = 16'h000a; // 0x3f8e
	13'h1fc8: q0 = 16'hee40; // 0x3f90
	13'h1fc9: q0 = 16'he640; // 0x3f92
	13'h1fca: q0 = 16'h3f00; // 0x3f94
	13'h1fcb: q0 = 16'h302e; // 0x3f96
	13'h1fcc: q0 = 16'h0008; // 0x3f98
	13'h1fcd: q0 = 16'hee40; // 0x3f9a
	13'h1fce: q0 = 16'he640; // 0x3f9c
	13'h1fcf: q0 = 16'h3f00; // 0x3f9e
	13'h1fd0: q0 = 16'h4eb9; // 0x3fa0
	13'h1fd1: q0 = 16'h0000; // 0x3fa2
	13'h1fd2: q0 = 16'h3d18; // 0x3fa4
	13'h1fd3: q0 = 16'h5c4f; // 0x3fa6
	13'h1fd4: q0 = 16'h4e5e; // 0x3fa8
	13'h1fd5: q0 = 16'h4e75; // 0x3faa
	13'h1fd6: q0 = 16'h4e56; // 0x3fac
	13'h1fd7: q0 = 16'hfffc; // 0x3fae
	13'h1fd8: q0 = 16'h0c79; // 0x3fb0
	13'h1fd9: q0 = 16'h0001; // 0x3fb2
	13'h1fda: q0 = 16'h0001; // 0x3fb4
	13'h1fdb: q0 = 16'h8678; // 0x3fb6
	13'h1fdc: q0 = 16'h6708; // 0x3fb8
	13'h1fdd: q0 = 16'h4a79; // 0x3fba
	13'h1fde: q0 = 16'h0001; // 0x3fbc
	13'h1fdf: q0 = 16'h867e; // 0x3fbe
	13'h1fe0: q0 = 16'h6604; // 0x3fc0
	13'h1fe1: q0 = 16'h7001; // 0x3fc2
	13'h1fe2: q0 = 16'h6002; // 0x3fc4
	13'h1fe3: q0 = 16'h4240; // 0x3fc6
	13'h1fe4: q0 = 16'h4e5e; // 0x3fc8
	13'h1fe5: q0 = 16'h4e75; // 0x3fca
	13'h1fe6: q0 = 16'h4e56; // 0x3fcc
	13'h1fe7: q0 = 16'h0000; // 0x3fce
	13'h1fe8: q0 = 16'h48e7; // 0x3fd0
	13'h1fe9: q0 = 16'h3f00; // 0x3fd2
	13'h1fea: q0 = 16'h3839; // 0x3fd4
	13'h1feb: q0 = 16'h0001; // 0x3fd6
	13'h1fec: q0 = 16'h81fc; // 0x3fd8
	13'h1fed: q0 = 16'h3c39; // 0x3fda
	13'h1fee: q0 = 16'h0001; // 0x3fdc
	13'h1fef: q0 = 16'h8936; // 0x3fde
	13'h1ff0: q0 = 16'h3a39; // 0x3fe0
	13'h1ff1: q0 = 16'h0001; // 0x3fe2
	13'h1ff2: q0 = 16'h8938; // 0x3fe4
	13'h1ff3: q0 = 16'h3e04; // 0x3fe6
	13'h1ff4: q0 = 16'he447; // 0x3fe8
	13'h1ff5: q0 = 16'h5247; // 0x3fea
	13'h1ff6: q0 = 16'hbe7c; // 0x3fec
	13'h1ff7: q0 = 16'h0008; // 0x3fee
	13'h1ff8: q0 = 16'h6f02; // 0x3ff0
	13'h1ff9: q0 = 16'h7e08; // 0x3ff2
	13'h1ffa: q0 = 16'h4a44; // 0x3ff4
	13'h1ffb: q0 = 16'h6602; // 0x3ff6
	13'h1ffc: q0 = 16'h4247; // 0x3ff8
	13'h1ffd: q0 = 16'h4eb9; // 0x3ffa
	13'h1ffe: q0 = 16'h0000; // 0x3ffc
	13'h1fff: q0 = 16'h4ec6; // 0x3ffe
  endcase

  always @(posedge clk)
    case (a)
	// foodfight code 136020-204.9d, 136020-303.8d
	13'h0000: q1 = 16'hb07c; // 0x0000
	13'h0001: q1 = 16'h0005; // 0x0002
	13'h0002: q1 = 16'h6732; // 0x0004
	13'h0003: q1 = 16'h3ebc; // 0x0006
	13'h0004: q1 = 16'h0020; // 0x0008
	13'h0005: q1 = 16'h3007; // 0x000a
	13'h0006: q1 = 16'he340; // 0x000c
	13'h0007: q1 = 16'h48c0; // 0x000e
	13'h0008: q1 = 16'h2f00; // 0x0010
	13'h0009: q1 = 16'h2039; // 0x0012
	13'h000a: q1 = 16'h0001; // 0x0014
	13'h000b: q1 = 16'h7f24; // 0x0016
	13'h000c: q1 = 16'hd0bc; // 0x0018
	13'h000d: q1 = 16'h0000; // 0x001a
	13'h000e: q1 = 16'h0012; // 0x001c
	13'h000f: q1 = 16'h5580; // 0x001e
	13'h0010: q1 = 16'h221f; // 0x0020
	13'h0011: q1 = 16'h9081; // 0x0022
	13'h0012: q1 = 16'h2040; // 0x0024
	13'h0013: q1 = 16'h3f10; // 0x0026
	13'h0014: q1 = 16'h3f05; // 0x0028
	13'h0015: q1 = 16'h0657; // 0x002a
	13'h0016: q1 = 16'h0400; // 0x002c
	13'h0017: q1 = 16'h3f06; // 0x002e
	13'h0018: q1 = 16'h4eb9; // 0x0030
	13'h0019: q1 = 16'h0000; // 0x0032
	13'h001a: q1 = 16'h3f80; // 0x0034
	13'h001b: q1 = 16'h5c4f; // 0x0036
	13'h001c: q1 = 16'hb87c; // 0x0038
	13'h001d: q1 = 16'h0008; // 0x003a
	13'h001e: q1 = 16'h6628; // 0x003c
	13'h001f: q1 = 16'h4a79; // 0x003e
	13'h0020: q1 = 16'h0001; // 0x0040
	13'h0021: q1 = 16'h81f4; // 0x0042
	13'h0022: q1 = 16'h6620; // 0x0044
	13'h0023: q1 = 16'h4eb9; // 0x0046
	13'h0024: q1 = 16'h0000; // 0x0048
	13'h0025: q1 = 16'h4ec6; // 0x004a
	13'h0026: q1 = 16'hb07c; // 0x004c
	13'h0027: q1 = 16'h0005; // 0x004e
	13'h0028: q1 = 16'h6714; // 0x0050
	13'h0029: q1 = 16'h2ebc; // 0x0052
	13'h002a: q1 = 16'h0000; // 0x0054
	13'h002b: q1 = 16'hc15a; // 0x0056
	13'h002c: q1 = 16'h4eb9; // 0x0058
	13'h002d: q1 = 16'h0000; // 0x005a
	13'h002e: q1 = 16'h7ff8; // 0x005c
	13'h002f: q1 = 16'h33fc; // 0x005e
	13'h0030: q1 = 16'h0001; // 0x0060
	13'h0031: q1 = 16'h0001; // 0x0062
	13'h0032: q1 = 16'h81f4; // 0x0064
	13'h0033: q1 = 16'h4a79; // 0x0066
	13'h0034: q1 = 16'h0001; // 0x0068
	13'h0035: q1 = 16'h867e; // 0x006a
	13'h0036: q1 = 16'h6652; // 0x006c
	13'h0037: q1 = 16'h4a44; // 0x006e
	13'h0038: q1 = 16'h664e; // 0x0070
	13'h0039: q1 = 16'h4eb9; // 0x0072
	13'h003a: q1 = 16'h0000; // 0x0074
	13'h003b: q1 = 16'h4ec6; // 0x0076
	13'h003c: q1 = 16'hb07c; // 0x0078
	13'h003d: q1 = 16'h0005; // 0x007a
	13'h003e: q1 = 16'h6742; // 0x007c
	13'h003f: q1 = 16'h4a79; // 0x007e
	13'h0040: q1 = 16'h0001; // 0x0080
	13'h0041: q1 = 16'h8058; // 0x0082
	13'h0042: q1 = 16'h6608; // 0x0084
	13'h0043: q1 = 16'h33fc; // 0x0086
	13'h0044: q1 = 16'h000f; // 0x0088
	13'h0045: q1 = 16'h0001; // 0x008a
	13'h0046: q1 = 16'h8058; // 0x008c
	13'h0047: q1 = 16'h5379; // 0x008e
	13'h0048: q1 = 16'h0001; // 0x0090
	13'h0049: q1 = 16'h8058; // 0x0092
	13'h004a: q1 = 16'h0c79; // 0x0094
	13'h004b: q1 = 16'h0007; // 0x0096
	13'h004c: q1 = 16'h0001; // 0x0098
	13'h004d: q1 = 16'h8058; // 0x009a
	13'h004e: q1 = 16'h6c06; // 0x009c
	13'h004f: q1 = 16'h363c; // 0x009e
	13'h0050: q1 = 16'h008a; // 0x00a0
	13'h0051: q1 = 16'h6002; // 0x00a2
	13'h0052: q1 = 16'h7640; // 0x00a4
	13'h0053: q1 = 16'h3ebc; // 0x00a6
	13'h0054: q1 = 16'h003e; // 0x00a8
	13'h0055: q1 = 16'h3f03; // 0x00aa
	13'h0056: q1 = 16'h3f05; // 0x00ac
	13'h0057: q1 = 16'h0657; // 0x00ae
	13'h0058: q1 = 16'h0400; // 0x00b0
	13'h0059: q1 = 16'h3f06; // 0x00b2
	13'h005a: q1 = 16'h4eb9; // 0x00b4
	13'h005b: q1 = 16'h0000; // 0x00b6
	13'h005c: q1 = 16'h3f80; // 0x00b8
	13'h005d: q1 = 16'h5c4f; // 0x00ba
	13'h005e: q1 = 16'h6000; // 0x00bc
	13'h005f: q1 = 16'h009a; // 0x00be
	13'h0060: q1 = 16'h0c79; // 0x00c0
	13'h0061: q1 = 16'h0001; // 0x00c2
	13'h0062: q1 = 16'h0001; // 0x00c4
	13'h0063: q1 = 16'h8678; // 0x00c6
	13'h0064: q1 = 16'h6700; // 0x00c8
	13'h0065: q1 = 16'h008e; // 0x00ca
	13'h0066: q1 = 16'h4a79; // 0x00cc
	13'h0067: q1 = 16'h0001; // 0x00ce
	13'h0068: q1 = 16'h8058; // 0x00d0
	13'h0069: q1 = 16'h666a; // 0x00d2
	13'h006a: q1 = 16'h5279; // 0x00d4
	13'h006b: q1 = 16'h0001; // 0x00d6
	13'h006c: q1 = 16'h867e; // 0x00d8
	13'h006d: q1 = 16'h0c79; // 0x00da
	13'h006e: q1 = 16'h000a; // 0x00dc
	13'h006f: q1 = 16'h0001; // 0x00de
	13'h0070: q1 = 16'h867e; // 0x00e0
	13'h0071: q1 = 16'h6f06; // 0x00e2
	13'h0072: q1 = 16'h4279; // 0x00e4
	13'h0073: q1 = 16'h0001; // 0x00e6
	13'h0074: q1 = 16'h867e; // 0x00e8
	13'h0075: q1 = 16'h3039; // 0x00ea
	13'h0076: q1 = 16'h0001; // 0x00ec
	13'h0077: q1 = 16'h867e; // 0x00ee
	13'h0078: q1 = 16'he340; // 0x00f0
	13'h0079: q1 = 16'h48c0; // 0x00f2
	13'h007a: q1 = 16'hd0bc; // 0x00f4
	13'h007b: q1 = 16'h0000; // 0x00f6
	13'h007c: q1 = 16'hcab2; // 0x00f8
	13'h007d: q1 = 16'h2040; // 0x00fa
	13'h007e: q1 = 16'h33d0; // 0x00fc
	13'h007f: q1 = 16'h0001; // 0x00fe
	13'h0080: q1 = 16'h8058; // 0x0100
	13'h0081: q1 = 16'h0c79; // 0x0102
	13'h0082: q1 = 16'h0009; // 0x0104
	13'h0083: q1 = 16'h0001; // 0x0106
	13'h0084: q1 = 16'h867e; // 0x0108
	13'h0085: q1 = 16'h660c; // 0x010a
	13'h0086: q1 = 16'h2ebc; // 0x010c
	13'h0087: q1 = 16'h0000; // 0x010e
	13'h0088: q1 = 16'hc7bc; // 0x0110
	13'h0089: q1 = 16'h4eb9; // 0x0112
	13'h008a: q1 = 16'h0000; // 0x0114
	13'h008b: q1 = 16'h7dd8; // 0x0116
	13'h008c: q1 = 16'h3ebc; // 0x0118
	13'h008d: q1 = 16'h0021; // 0x011a
	13'h008e: q1 = 16'h3039; // 0x011c
	13'h008f: q1 = 16'h0001; // 0x011e
	13'h0090: q1 = 16'h867e; // 0x0120
	13'h0091: q1 = 16'he340; // 0x0122
	13'h0092: q1 = 16'h48c0; // 0x0124
	13'h0093: q1 = 16'hd0bc; // 0x0126
	13'h0094: q1 = 16'h0000; // 0x0128
	13'h0095: q1 = 16'hca9c; // 0x012a
	13'h0096: q1 = 16'h2040; // 0x012c
	13'h0097: q1 = 16'h3f10; // 0x012e
	13'h0098: q1 = 16'h3f05; // 0x0130
	13'h0099: q1 = 16'h3f06; // 0x0132
	13'h009a: q1 = 16'h4eb9; // 0x0134
	13'h009b: q1 = 16'h0000; // 0x0136
	13'h009c: q1 = 16'h3f80; // 0x0138
	13'h009d: q1 = 16'h5c4f; // 0x013a
	13'h009e: q1 = 16'h6006; // 0x013c
	13'h009f: q1 = 16'h5379; // 0x013e
	13'h00a0: q1 = 16'h0001; // 0x0140
	13'h00a1: q1 = 16'h8058; // 0x0142
	13'h00a2: q1 = 16'h4a44; // 0x0144
	13'h00a3: q1 = 16'h6610; // 0x0146
	13'h00a4: q1 = 16'h4a79; // 0x0148
	13'h00a5: q1 = 16'h0001; // 0x014a
	13'h00a6: q1 = 16'h867e; // 0x014c
	13'h00a7: q1 = 16'h6608; // 0x014e
	13'h00a8: q1 = 16'h33fc; // 0x0150
	13'h00a9: q1 = 16'h000f; // 0x0152
	13'h00aa: q1 = 16'h0001; // 0x0154
	13'h00ab: q1 = 16'h8058; // 0x0156
	13'h00ac: q1 = 16'h4a9f; // 0x0158
	13'h00ad: q1 = 16'h4cdf; // 0x015a
	13'h00ae: q1 = 16'h00f8; // 0x015c
	13'h00af: q1 = 16'h4e5e; // 0x015e
	13'h00b0: q1 = 16'h4e75; // 0x0160
	13'h00b1: q1 = 16'h4e56; // 0x0162
	13'h00b2: q1 = 16'hfffc; // 0x0164
	13'h00b3: q1 = 16'h3ebc; // 0x0166
	13'h00b4: q1 = 16'h0001; // 0x0168
	13'h00b5: q1 = 16'h3f3c; // 0x016a
	13'h00b6: q1 = 16'h0040; // 0x016c
	13'h00b7: q1 = 16'h3f39; // 0x016e
	13'h00b8: q1 = 16'h0001; // 0x0170
	13'h00b9: q1 = 16'h8938; // 0x0172
	13'h00ba: q1 = 16'h0657; // 0x0174
	13'h00bb: q1 = 16'h0400; // 0x0176
	13'h00bc: q1 = 16'h3f39; // 0x0178
	13'h00bd: q1 = 16'h0001; // 0x017a
	13'h00be: q1 = 16'h8936; // 0x017c
	13'h00bf: q1 = 16'h4eb9; // 0x017e
	13'h00c0: q1 = 16'h0000; // 0x0180
	13'h00c1: q1 = 16'h3f80; // 0x0182
	13'h00c2: q1 = 16'h5c4f; // 0x0184
	13'h00c3: q1 = 16'h3ebc; // 0x0186
	13'h00c4: q1 = 16'h0001; // 0x0188
	13'h00c5: q1 = 16'h3f3c; // 0x018a
	13'h00c6: q1 = 16'h0040; // 0x018c
	13'h00c7: q1 = 16'h3f39; // 0x018e
	13'h00c8: q1 = 16'h0001; // 0x0190
	13'h00c9: q1 = 16'h8938; // 0x0192
	13'h00ca: q1 = 16'h3f39; // 0x0194
	13'h00cb: q1 = 16'h0001; // 0x0196
	13'h00cc: q1 = 16'h8936; // 0x0198
	13'h00cd: q1 = 16'h4eb9; // 0x019a
	13'h00ce: q1 = 16'h0000; // 0x019c
	13'h00cf: q1 = 16'h3f80; // 0x019e
	13'h00d0: q1 = 16'h5c4f; // 0x01a0
	13'h00d1: q1 = 16'h33fc; // 0x01a2
	13'h00d2: q1 = 16'h0001; // 0x01a4
	13'h00d3: q1 = 16'h0001; // 0x01a6
	13'h00d4: q1 = 16'h8678; // 0x01a8
	13'h00d5: q1 = 16'h4e5e; // 0x01aa
	13'h00d6: q1 = 16'h4e75; // 0x01ac
	13'h00d7: q1 = 16'h4e56; // 0x01ae
	13'h00d8: q1 = 16'hfff8; // 0x01b0
	13'h00d9: q1 = 16'h48e7; // 0x01b2
	13'h00da: q1 = 16'h0104; // 0x01b4
	13'h00db: q1 = 16'h2a79; // 0x01b6
	13'h00dc: q1 = 16'h0001; // 0x01b8
	13'h00dd: q1 = 16'h7fb8; // 0x01ba
	13'h00de: q1 = 16'h33fc; // 0x01bc
	13'h00df: q1 = 16'h0580; // 0x01be
	13'h00e0: q1 = 16'h0001; // 0x01c0
	13'h00e1: q1 = 16'h8936; // 0x01c2
	13'h00e2: q1 = 16'h0c55; // 0x01c4
	13'h00e3: q1 = 16'h0006; // 0x01c6
	13'h00e4: q1 = 16'h6f1c; // 0x01c8
	13'h00e5: q1 = 16'h3ebc; // 0x01ca
	13'h00e6: q1 = 16'h7000; // 0x01cc
	13'h00e7: q1 = 16'h3f3c; // 0x01ce
	13'h00e8: q1 = 16'h1400; // 0x01d0
	13'h00e9: q1 = 16'h4eb9; // 0x01d2
	13'h00ea: q1 = 16'h0000; // 0x01d4
	13'h00eb: q1 = 16'h8e6c; // 0x01d6
	13'h00ec: q1 = 16'h4a5f; // 0x01d8
	13'h00ed: q1 = 16'hd07c; // 0x01da
	13'h00ee: q1 = 16'h0400; // 0x01dc
	13'h00ef: q1 = 16'h33c0; // 0x01de
	13'h00f0: q1 = 16'h0001; // 0x01e0
	13'h00f1: q1 = 16'h8938; // 0x01e2
	13'h00f2: q1 = 16'h6008; // 0x01e4
	13'h00f3: q1 = 16'h33fc; // 0x01e6
	13'h00f4: q1 = 16'h4400; // 0x01e8
	13'h00f5: q1 = 16'h0001; // 0x01ea
	13'h00f6: q1 = 16'h8938; // 0x01ec
	13'h00f7: q1 = 16'h2ebc; // 0x01ee
	13'h00f8: q1 = 16'h0001; // 0x01f0
	13'h00f9: q1 = 16'h8938; // 0x01f2
	13'h00fa: q1 = 16'h2f3c; // 0x01f4
	13'h00fb: q1 = 16'h0001; // 0x01f6
	13'h00fc: q1 = 16'h8936; // 0x01f8
	13'h00fd: q1 = 16'h4eb9; // 0x01fa
	13'h00fe: q1 = 16'h0000; // 0x01fc
	13'h00ff: q1 = 16'hbee0; // 0x01fe
	13'h0100: q1 = 16'h4a9f; // 0x0200
	13'h0101: q1 = 16'h3ebc; // 0x0202
	13'h0102: q1 = 16'h0020; // 0x0204
	13'h0103: q1 = 16'h200e; // 0x0206
	13'h0104: q1 = 16'hd0bc; // 0x0208
	13'h0105: q1 = 16'hffff; // 0x020a
	13'h0106: q1 = 16'hfff8; // 0x020c
	13'h0107: q1 = 16'h2f00; // 0x020e
	13'h0108: q1 = 16'h200e; // 0x0210
	13'h0109: q1 = 16'hd0bc; // 0x0212
	13'h010a: q1 = 16'hffff; // 0x0214
	13'h010b: q1 = 16'hfffe; // 0x0216
	13'h010c: q1 = 16'h2f00; // 0x0218
	13'h010d: q1 = 16'h3f15; // 0x021a
	13'h010e: q1 = 16'h4eb9; // 0x021c
	13'h010f: q1 = 16'h0000; // 0x021e
	13'h0110: q1 = 16'h1402; // 0x0220
	13'h0111: q1 = 16'hdefc; // 0x0222
	13'h0112: q1 = 16'h000a; // 0x0224
	13'h0113: q1 = 16'h302e; // 0x0226
	13'h0114: q1 = 16'hfffe; // 0x0228
	13'h0115: q1 = 16'h5340; // 0x022a
	13'h0116: q1 = 16'hc1fc; // 0x022c
	13'h0117: q1 = 16'h0012; // 0x022e
	13'h0118: q1 = 16'hd0bc; // 0x0230
	13'h0119: q1 = 16'h0000; // 0x0232
	13'h011a: q1 = 16'hcac8; // 0x0234
	13'h011b: q1 = 16'h23c0; // 0x0236
	13'h011c: q1 = 16'h0001; // 0x0238
	13'h011d: q1 = 16'h7f24; // 0x023a
	13'h011e: q1 = 16'h33ee; // 0x023c
	13'h011f: q1 = 16'hfff8; // 0x023e
	13'h0120: q1 = 16'h0001; // 0x0240
	13'h0121: q1 = 16'h76f2; // 0x0242
	13'h0122: q1 = 16'h3e95; // 0x0244
	13'h0123: q1 = 16'h4eb9; // 0x0246
	13'h0124: q1 = 16'h0000; // 0x0248
	13'h0125: q1 = 16'h14d0; // 0x024a
	13'h0126: q1 = 16'h4279; // 0x024c
	13'h0127: q1 = 16'h0001; // 0x024e
	13'h0128: q1 = 16'h8678; // 0x0250
	13'h0129: q1 = 16'h4279; // 0x0252
	13'h012a: q1 = 16'h0001; // 0x0254
	13'h012b: q1 = 16'h81f4; // 0x0256
	13'h012c: q1 = 16'h33fc; // 0x0258
	13'h012d: q1 = 16'h0001; // 0x025a
	13'h012e: q1 = 16'h0001; // 0x025c
	13'h012f: q1 = 16'h8a78; // 0x025e
	13'h0130: q1 = 16'h4279; // 0x0260
	13'h0131: q1 = 16'h0001; // 0x0262
	13'h0132: q1 = 16'h867e; // 0x0264
	13'h0133: q1 = 16'h33f9; // 0x0266
	13'h0134: q1 = 16'h0000; // 0x0268
	13'h0135: q1 = 16'hcab2; // 0x026a
	13'h0136: q1 = 16'h0001; // 0x026c
	13'h0137: q1 = 16'h8058; // 0x026e
	13'h0138: q1 = 16'h3ebc; // 0x0270
	13'h0139: q1 = 16'h0021; // 0x0272
	13'h013a: q1 = 16'h3f39; // 0x0274
	13'h013b: q1 = 16'h0000; // 0x0276
	13'h013c: q1 = 16'hca9c; // 0x0278
	13'h013d: q1 = 16'h3f39; // 0x027a
	13'h013e: q1 = 16'h0001; // 0x027c
	13'h013f: q1 = 16'h8938; // 0x027e
	13'h0140: q1 = 16'h3f39; // 0x0280
	13'h0141: q1 = 16'h0001; // 0x0282
	13'h0142: q1 = 16'h8936; // 0x0284
	13'h0143: q1 = 16'h4eb9; // 0x0286
	13'h0144: q1 = 16'h0000; // 0x0288
	13'h0145: q1 = 16'h3f80; // 0x028a
	13'h0146: q1 = 16'h5c4f; // 0x028c
	13'h0147: q1 = 16'h3ebc; // 0x028e
	13'h0148: q1 = 16'h0020; // 0x0290
	13'h0149: q1 = 16'h2079; // 0x0292
	13'h014a: q1 = 16'h0001; // 0x0294
	13'h014b: q1 = 16'h7f24; // 0x0296
	13'h014c: q1 = 16'h3f10; // 0x0298
	13'h014d: q1 = 16'h3f39; // 0x029a
	13'h014e: q1 = 16'h0001; // 0x029c
	13'h014f: q1 = 16'h8938; // 0x029e
	13'h0150: q1 = 16'h0657; // 0x02a0
	13'h0151: q1 = 16'h0400; // 0x02a2
	13'h0152: q1 = 16'h3f39; // 0x02a4
	13'h0153: q1 = 16'h0001; // 0x02a6
	13'h0154: q1 = 16'h8936; // 0x02a8
	13'h0155: q1 = 16'h4eb9; // 0x02aa
	13'h0156: q1 = 16'h0000; // 0x02ac
	13'h0157: q1 = 16'h3f80; // 0x02ae
	13'h0158: q1 = 16'h5c4f; // 0x02b0
	13'h0159: q1 = 16'h4a9f; // 0x02b2
	13'h015a: q1 = 16'h4cdf; // 0x02b4
	13'h015b: q1 = 16'h2000; // 0x02b6
	13'h015c: q1 = 16'h4e5e; // 0x02b8
	13'h015d: q1 = 16'h4e75; // 0x02ba
	13'h015e: q1 = 16'h4e56; // 0x02bc
	13'h015f: q1 = 16'hfffc; // 0x02be
	13'h0160: q1 = 16'h33fc; // 0x02c0
	13'h0161: q1 = 16'h0580; // 0x02c2
	13'h0162: q1 = 16'h0001; // 0x02c4
	13'h0163: q1 = 16'h8936; // 0x02c6
	13'h0164: q1 = 16'h33fc; // 0x02c8
	13'h0165: q1 = 16'h4400; // 0x02ca
	13'h0166: q1 = 16'h0001; // 0x02cc
	13'h0167: q1 = 16'h8938; // 0x02ce
	13'h0168: q1 = 16'h4e5e; // 0x02d0
	13'h0169: q1 = 16'h4e75; // 0x02d2
	13'h016a: q1 = 16'h4e56; // 0x02d4
	13'h016b: q1 = 16'h0000; // 0x02d6
	13'h016c: q1 = 16'h48e7; // 0x02d8
	13'h016d: q1 = 16'h0700; // 0x02da
	13'h016e: q1 = 16'h3e2e; // 0x02dc
	13'h016f: q1 = 16'h0008; // 0x02de
	13'h0170: q1 = 16'h9e79; // 0x02e0
	13'h0171: q1 = 16'h0001; // 0x02e2
	13'h0172: q1 = 16'h8936; // 0x02e4
	13'h0173: q1 = 16'h4a47; // 0x02e6
	13'h0174: q1 = 16'h6c06; // 0x02e8
	13'h0175: q1 = 16'h3007; // 0x02ea
	13'h0176: q1 = 16'h4440; // 0x02ec
	13'h0177: q1 = 16'h3e00; // 0x02ee
	13'h0178: q1 = 16'h4a6e; // 0x02f0
	13'h0179: q1 = 16'h000c; // 0x02f2
	13'h017a: q1 = 16'h6706; // 0x02f4
	13'h017b: q1 = 16'h3c3c; // 0x02f6
	13'h017c: q1 = 16'h1000; // 0x02f8
	13'h017d: q1 = 16'h6004; // 0x02fa
	13'h017e: q1 = 16'h3c3c; // 0x02fc
	13'h017f: q1 = 16'h0400; // 0x02fe
	13'h0180: q1 = 16'hbe46; // 0x0300
	13'h0181: q1 = 16'h6f04; // 0x0302
	13'h0182: q1 = 16'h4240; // 0x0304
	13'h0183: q1 = 16'h602e; // 0x0306
	13'h0184: q1 = 16'h3e2e; // 0x0308
	13'h0185: q1 = 16'h000a; // 0x030a
	13'h0186: q1 = 16'h9e79; // 0x030c
	13'h0187: q1 = 16'h0001; // 0x030e
	13'h0188: q1 = 16'h8938; // 0x0310
	13'h0189: q1 = 16'h4a47; // 0x0312
	13'h018a: q1 = 16'h6c06; // 0x0314
	13'h018b: q1 = 16'h3007; // 0x0316
	13'h018c: q1 = 16'h4440; // 0x0318
	13'h018d: q1 = 16'h3e00; // 0x031a
	13'h018e: q1 = 16'h4a6e; // 0x031c
	13'h018f: q1 = 16'h000c; // 0x031e
	13'h0190: q1 = 16'h6706; // 0x0320
	13'h0191: q1 = 16'h3c3c; // 0x0322
	13'h0192: q1 = 16'h1000; // 0x0324
	13'h0193: q1 = 16'h6004; // 0x0326
	13'h0194: q1 = 16'h3c3c; // 0x0328
	13'h0195: q1 = 16'h0600; // 0x032a
	13'h0196: q1 = 16'hbe46; // 0x032c
	13'h0197: q1 = 16'h6f04; // 0x032e
	13'h0198: q1 = 16'h4240; // 0x0330
	13'h0199: q1 = 16'h6002; // 0x0332
	13'h019a: q1 = 16'h7001; // 0x0334
	13'h019b: q1 = 16'h4a9f; // 0x0336
	13'h019c: q1 = 16'h4cdf; // 0x0338
	13'h019d: q1 = 16'h00c0; // 0x033a
	13'h019e: q1 = 16'h4e5e; // 0x033c
	13'h019f: q1 = 16'h4e75; // 0x033e
	13'h01a0: q1 = 16'h4e56; // 0x0340
	13'h01a1: q1 = 16'hfffa; // 0x0342
	13'h01a2: q1 = 16'h48e7; // 0x0344
	13'h01a3: q1 = 16'h0704; // 0x0346
	13'h01a4: q1 = 16'h4a79; // 0x0348
	13'h01a5: q1 = 16'h0001; // 0x034a
	13'h01a6: q1 = 16'h8676; // 0x034c
	13'h01a7: q1 = 16'h6600; // 0x034e
	13'h01a8: q1 = 16'h00ec; // 0x0350
	13'h01a9: q1 = 16'h2079; // 0x0352
	13'h01aa: q1 = 16'h0001; // 0x0354
	13'h01ab: q1 = 16'h7fb8; // 0x0356
	13'h01ac: q1 = 16'h3010; // 0x0358
	13'h01ad: q1 = 16'he540; // 0x035a
	13'h01ae: q1 = 16'h2279; // 0x035c
	13'h01af: q1 = 16'h0001; // 0x035e
	13'h01b0: q1 = 16'h7fb8; // 0x0360
	13'h01b1: q1 = 16'hd051; // 0x0362
	13'h01b2: q1 = 16'h3c00; // 0x0364
	13'h01b3: q1 = 16'hbc7c; // 0x0366
	13'h01b4: q1 = 16'h00fa; // 0x0368
	13'h01b5: q1 = 16'h6f04; // 0x036a
	13'h01b6: q1 = 16'h3c3c; // 0x036c
	13'h01b7: q1 = 16'h00fa; // 0x036e
	13'h01b8: q1 = 16'h200e; // 0x0370
	13'h01b9: q1 = 16'hd0bc; // 0x0372
	13'h01ba: q1 = 16'hffff; // 0x0374
	13'h01bb: q1 = 16'hfffa; // 0x0376
	13'h01bc: q1 = 16'h2e80; // 0x0378
	13'h01bd: q1 = 16'h3f06; // 0x037a
	13'h01be: q1 = 16'h4eb9; // 0x037c
	13'h01bf: q1 = 16'h0000; // 0x037e
	13'h01c0: q1 = 16'h0828; // 0x0380
	13'h01c1: q1 = 16'h4a5f; // 0x0382
	13'h01c2: q1 = 16'h2ebc; // 0x0384
	13'h01c3: q1 = 16'h0000; // 0x0386
	13'h01c4: q1 = 16'hca0c; // 0x0388
	13'h01c5: q1 = 16'h200e; // 0x038a
	13'h01c6: q1 = 16'hd0bc; // 0x038c
	13'h01c7: q1 = 16'hffff; // 0x038e
	13'h01c8: q1 = 16'hfffa; // 0x0390
	13'h01c9: q1 = 16'h2f00; // 0x0392
	13'h01ca: q1 = 16'h4eb9; // 0x0394
	13'h01cb: q1 = 16'h0000; // 0x0396
	13'h01cc: q1 = 16'h0770; // 0x0398
	13'h01cd: q1 = 16'h4a9f; // 0x039a
	13'h01ce: q1 = 16'h4a79; // 0x039c
	13'h01cf: q1 = 16'h0001; // 0x039e
	13'h01d0: q1 = 16'h8a78; // 0x03a0
	13'h01d1: q1 = 16'h6750; // 0x03a2
	13'h01d2: q1 = 16'h4247; // 0x03a4
	13'h01d3: q1 = 16'hbe7c; // 0x03a6
	13'h01d4: q1 = 16'h0005; // 0x03a8
	13'h01d5: q1 = 16'h6c48; // 0x03aa
	13'h01d6: q1 = 16'h3007; // 0x03ac
	13'h01d7: q1 = 16'he340; // 0x03ae
	13'h01d8: q1 = 16'h48c0; // 0x03b0
	13'h01d9: q1 = 16'hd0bc; // 0x03b2
	13'h01da: q1 = 16'h0001; // 0x03b4
	13'h01db: q1 = 16'h8694; // 0x03b6
	13'h01dc: q1 = 16'h2e80; // 0x03b8
	13'h01dd: q1 = 16'h3007; // 0x03ba
	13'h01de: q1 = 16'he340; // 0x03bc
	13'h01df: q1 = 16'h48c0; // 0x03be
	13'h01e0: q1 = 16'hd0bc; // 0x03c0
	13'h01e1: q1 = 16'h0001; // 0x03c2
	13'h01e2: q1 = 16'h869e; // 0x03c4
	13'h01e3: q1 = 16'h2f00; // 0x03c6
	13'h01e4: q1 = 16'h3f39; // 0x03c8
	13'h01e5: q1 = 16'h0001; // 0x03ca
	13'h01e6: q1 = 16'h8938; // 0x03cc
	13'h01e7: q1 = 16'h0657; // 0x03ce
	13'h01e8: q1 = 16'h0400; // 0x03d0
	13'h01e9: q1 = 16'h3007; // 0x03d2
	13'h01ea: q1 = 16'h4281; // 0x03d4
	13'h01eb: q1 = 16'h720a; // 0x03d6
	13'h01ec: q1 = 16'he360; // 0x03d8
	13'h01ed: q1 = 16'h3f00; // 0x03da
	13'h01ee: q1 = 16'h3039; // 0x03dc
	13'h01ef: q1 = 16'h0001; // 0x03de
	13'h01f0: q1 = 16'h8936; // 0x03e0
	13'h01f1: q1 = 16'hd157; // 0x03e2
	13'h01f2: q1 = 16'h0657; // 0x03e4
	13'h01f3: q1 = 16'h0800; // 0x03e6
	13'h01f4: q1 = 16'h4eb9; // 0x03e8
	13'h01f5: q1 = 16'h0000; // 0x03ea
	13'h01f6: q1 = 16'h3dbe; // 0x03ec
	13'h01f7: q1 = 16'hbf8f; // 0x03ee
	13'h01f8: q1 = 16'h5247; // 0x03f0
	13'h01f9: q1 = 16'h60b2; // 0x03f2
	13'h01fa: q1 = 16'h4279; // 0x03f4
	13'h01fb: q1 = 16'h0001; // 0x03f6
	13'h01fc: q1 = 16'h8a78; // 0x03f8
	13'h01fd: q1 = 16'h4247; // 0x03fa
	13'h01fe: q1 = 16'h4bee; // 0x03fc
	13'h01ff: q1 = 16'hfffa; // 0x03fe
	13'h0200: q1 = 16'h4a15; // 0x0400
	13'h0201: q1 = 16'h6738; // 0x0402
	13'h0202: q1 = 16'h1c15; // 0x0404
	13'h0203: q1 = 16'h4886; // 0x0406
	13'h0204: q1 = 16'h3ebc; // 0x0408
	13'h0205: q1 = 16'h0036; // 0x040a
	13'h0206: q1 = 16'h3f06; // 0x040c
	13'h0207: q1 = 16'h3f39; // 0x040e
	13'h0208: q1 = 16'h0001; // 0x0410
	13'h0209: q1 = 16'h8938; // 0x0412
	13'h020a: q1 = 16'h0657; // 0x0414
	13'h020b: q1 = 16'h0400; // 0x0416
	13'h020c: q1 = 16'h3007; // 0x0418
	13'h020d: q1 = 16'h4281; // 0x041a
	13'h020e: q1 = 16'h720a; // 0x041c
	13'h020f: q1 = 16'he360; // 0x041e
	13'h0210: q1 = 16'h3f00; // 0x0420
	13'h0211: q1 = 16'h3039; // 0x0422
	13'h0212: q1 = 16'h0001; // 0x0424
	13'h0213: q1 = 16'h8936; // 0x0426
	13'h0214: q1 = 16'hd157; // 0x0428
	13'h0215: q1 = 16'h0657; // 0x042a
	13'h0216: q1 = 16'h0800; // 0x042c
	13'h0217: q1 = 16'h4eb9; // 0x042e
	13'h0218: q1 = 16'h0000; // 0x0430
	13'h0219: q1 = 16'h3f80; // 0x0432
	13'h021a: q1 = 16'h5c4f; // 0x0434
	13'h021b: q1 = 16'h5247; // 0x0436
	13'h021c: q1 = 16'h528d; // 0x0438
	13'h021d: q1 = 16'h60c4; // 0x043a
	13'h021e: q1 = 16'h4a9f; // 0x043c
	13'h021f: q1 = 16'h4cdf; // 0x043e
	13'h0220: q1 = 16'h20c0; // 0x0440
	13'h0221: q1 = 16'h4e5e; // 0x0442
	13'h0222: q1 = 16'h4e75; // 0x0444
	13'h0223: q1 = 16'h4e56; // 0x0446
	13'h0224: q1 = 16'h0000; // 0x0448
	13'h0225: q1 = 16'h48e7; // 0x044a
	13'h0226: q1 = 16'h0300; // 0x044c
	13'h0227: q1 = 16'h4247; // 0x044e
	13'h0228: q1 = 16'hbe7c; // 0x0450
	13'h0229: q1 = 16'h0005; // 0x0452
	13'h022a: q1 = 16'h6c4c; // 0x0454
	13'h022b: q1 = 16'h3007; // 0x0456
	13'h022c: q1 = 16'he340; // 0x0458
	13'h022d: q1 = 16'h48c0; // 0x045a
	13'h022e: q1 = 16'hd0bc; // 0x045c
	13'h022f: q1 = 16'h0001; // 0x045e
	13'h0230: q1 = 16'h8694; // 0x0460
	13'h0231: q1 = 16'h2040; // 0x0462
	13'h0232: q1 = 16'h3e90; // 0x0464
	13'h0233: q1 = 16'h3007; // 0x0466
	13'h0234: q1 = 16'he340; // 0x0468
	13'h0235: q1 = 16'h48c0; // 0x046a
	13'h0236: q1 = 16'hd0bc; // 0x046c
	13'h0237: q1 = 16'h0001; // 0x046e
	13'h0238: q1 = 16'h869e; // 0x0470
	13'h0239: q1 = 16'h2040; // 0x0472
	13'h023a: q1 = 16'h3f10; // 0x0474
	13'h023b: q1 = 16'h3f39; // 0x0476
	13'h023c: q1 = 16'h0001; // 0x0478
	13'h023d: q1 = 16'h8938; // 0x047a
	13'h023e: q1 = 16'h0657; // 0x047c
	13'h023f: q1 = 16'h0400; // 0x047e
	13'h0240: q1 = 16'h3007; // 0x0480
	13'h0241: q1 = 16'h4281; // 0x0482
	13'h0242: q1 = 16'h720a; // 0x0484
	13'h0243: q1 = 16'he360; // 0x0486
	13'h0244: q1 = 16'h3f00; // 0x0488
	13'h0245: q1 = 16'h3039; // 0x048a
	13'h0246: q1 = 16'h0001; // 0x048c
	13'h0247: q1 = 16'h8936; // 0x048e
	13'h0248: q1 = 16'hd157; // 0x0490
	13'h0249: q1 = 16'h0657; // 0x0492
	13'h024a: q1 = 16'h0800; // 0x0494
	13'h024b: q1 = 16'h4eb9; // 0x0496
	13'h024c: q1 = 16'h0000; // 0x0498
	13'h024d: q1 = 16'h3f80; // 0x049a
	13'h024e: q1 = 16'h5c4f; // 0x049c
	13'h024f: q1 = 16'h5247; // 0x049e
	13'h0250: q1 = 16'h60ae; // 0x04a0
	13'h0251: q1 = 16'h4a9f; // 0x04a2
	13'h0252: q1 = 16'h4cdf; // 0x04a4
	13'h0253: q1 = 16'h0080; // 0x04a6
	13'h0254: q1 = 16'h4e5e; // 0x04a8
	13'h0255: q1 = 16'h4e75; // 0x04aa
	13'h0256: q1 = 16'h4e56; // 0x04ac
	13'h0257: q1 = 16'hffe0; // 0x04ae
	13'h0258: q1 = 16'h48e7; // 0x04b0
	13'h0259: q1 = 16'h1f00; // 0x04b2
	13'h025a: q1 = 16'h0c79; // 0x04b4
	13'h025b: q1 = 16'h0002; // 0x04b6
	13'h025c: q1 = 16'h0001; // 0x04b8
	13'h025d: q1 = 16'h7f5e; // 0x04ba
	13'h025e: q1 = 16'h660a; // 0x04bc
	13'h025f: q1 = 16'h33fc; // 0x04be
	13'h0260: q1 = 16'h0002; // 0x04c0
	13'h0261: q1 = 16'h0001; // 0x04c2
	13'h0262: q1 = 16'h87dc; // 0x04c4
	13'h0263: q1 = 16'h6008; // 0x04c6
	13'h0264: q1 = 16'h33fc; // 0x04c8
	13'h0265: q1 = 16'h0001; // 0x04ca
	13'h0266: q1 = 16'h0001; // 0x04cc
	13'h0267: q1 = 16'h87dc; // 0x04ce
	13'h0268: q1 = 16'h4eb9; // 0x04d0
	13'h0269: q1 = 16'h0000; // 0x04d2
	13'h026a: q1 = 16'h1266; // 0x04d4
	13'h026b: q1 = 16'h4eb9; // 0x04d6
	13'h026c: q1 = 16'h0000; // 0x04d8
	13'h026d: q1 = 16'ha964; // 0x04da
	13'h026e: q1 = 16'h33f9; // 0x04dc
	13'h026f: q1 = 16'h0001; // 0x04de
	13'h0270: q1 = 16'h7eb6; // 0x04e0
	13'h0271: q1 = 16'h0001; // 0x04e2
	13'h0272: q1 = 16'h8628; // 0x04e4
	13'h0273: q1 = 16'h0c79; // 0x04e6
	13'h0274: q1 = 16'h0002; // 0x04e8
	13'h0275: q1 = 16'h0001; // 0x04ea
	13'h0276: q1 = 16'h87dc; // 0x04ec
	13'h0277: q1 = 16'h660a; // 0x04ee
	13'h0278: q1 = 16'h33f9; // 0x04f0
	13'h0279: q1 = 16'h0001; // 0x04f2
	13'h027a: q1 = 16'h7eb6; // 0x04f4
	13'h027b: q1 = 16'h0001; // 0x04f6
	13'h027c: q1 = 16'h864e; // 0x04f8
	13'h027d: q1 = 16'h0c79; // 0x04fa
	13'h027e: q1 = 16'h0001; // 0x04fc
	13'h027f: q1 = 16'h0001; // 0x04fe
	13'h0280: q1 = 16'h757c; // 0x0500
	13'h0281: q1 = 16'h6e06; // 0x0502
	13'h0282: q1 = 16'h4279; // 0x0504
	13'h0283: q1 = 16'h0001; // 0x0506
	13'h0284: q1 = 16'h757c; // 0x0508
	13'h0285: q1 = 16'h4eb9; // 0x050a
	13'h0286: q1 = 16'h0000; // 0x050c
	13'h0287: q1 = 16'h87c8; // 0x050e
	13'h0288: q1 = 16'h4eb9; // 0x0510
	13'h0289: q1 = 16'h0000; // 0x0512
	13'h028a: q1 = 16'h4754; // 0x0514
	13'h028b: q1 = 16'h4eb9; // 0x0516
	13'h028c: q1 = 16'h0000; // 0x0518
	13'h028d: q1 = 16'h33e6; // 0x051a
	13'h028e: q1 = 16'h4279; // 0x051c
	13'h028f: q1 = 16'h0001; // 0x051e
	13'h0290: q1 = 16'h8054; // 0x0520
	13'h0291: q1 = 16'h23fc; // 0x0522
	13'h0292: q1 = 16'h0001; // 0x0524
	13'h0293: q1 = 16'h8628; // 0x0526
	13'h0294: q1 = 16'h0001; // 0x0528
	13'h0295: q1 = 16'h7fb8; // 0x052a
	13'h0296: q1 = 16'h33fc; // 0x052c
	13'h0297: q1 = 16'h0001; // 0x052e
	13'h0298: q1 = 16'h0001; // 0x0530
	13'h0299: q1 = 16'h7fc8; // 0x0532
	13'h029a: q1 = 16'h33fc; // 0x0534
	13'h029b: q1 = 16'h0001; // 0x0536
	13'h029c: q1 = 16'h0001; // 0x0538
	13'h029d: q1 = 16'h7eb8; // 0x053a
	13'h029e: q1 = 16'h2079; // 0x053c
	13'h029f: q1 = 16'h0001; // 0x053e
	13'h02a0: q1 = 16'h7fb8; // 0x0540
	13'h02a1: q1 = 16'h4a68; // 0x0542
	13'h02a2: q1 = 16'h0022; // 0x0544
	13'h02a3: q1 = 16'h6710; // 0x0546
	13'h02a4: q1 = 16'h4eb9; // 0x0548
	13'h02a5: q1 = 16'h0000; // 0x054a
	13'h02a6: q1 = 16'h9570; // 0x054c
	13'h02a7: q1 = 16'h2079; // 0x054e
	13'h02a8: q1 = 16'h0001; // 0x0550
	13'h02a9: q1 = 16'h7fb8; // 0x0552
	13'h02aa: q1 = 16'h4268; // 0x0554
	13'h02ab: q1 = 16'h0022; // 0x0556
	13'h02ac: q1 = 16'h4eb9; // 0x0558
	13'h02ad: q1 = 16'h0000; // 0x055a
	13'h02ae: q1 = 16'h8ca4; // 0x055c
	13'h02af: q1 = 16'h2079; // 0x055e
	13'h02b0: q1 = 16'h0001; // 0x0560
	13'h02b1: q1 = 16'h7fb8; // 0x0562
	13'h02b2: q1 = 16'h5368; // 0x0564
	13'h02b3: q1 = 16'h0002; // 0x0566
	13'h02b4: q1 = 16'h2079; // 0x0568
	13'h02b5: q1 = 16'h0001; // 0x056a
	13'h02b6: q1 = 16'h7fb8; // 0x056c
	13'h02b7: q1 = 16'h4a68; // 0x056e
	13'h02b8: q1 = 16'h0002; // 0x0570
	13'h02b9: q1 = 16'h6600; // 0x0572
	13'h02ba: q1 = 16'h00e0; // 0x0574
	13'h02bb: q1 = 16'h4245; // 0x0576
	13'h02bc: q1 = 16'h783e; // 0x0578
	13'h02bd: q1 = 16'h2ebc; // 0x057a
	13'h02be: q1 = 16'h0000; // 0x057c
	13'h02bf: q1 = 16'hcedc; // 0x057e
	13'h02c0: q1 = 16'h4eb9; // 0x0580
	13'h02c1: q1 = 16'h0000; // 0x0582
	13'h02c2: q1 = 16'h7ff8; // 0x0584
	13'h02c3: q1 = 16'h3ebc; // 0x0586
	13'h02c4: q1 = 16'h002e; // 0x0588
	13'h02c5: q1 = 16'h200e; // 0x058a
	13'h02c6: q1 = 16'hd0bc; // 0x058c
	13'h02c7: q1 = 16'hffff; // 0x058e
	13'h02c8: q1 = 16'hffe0; // 0x0590
	13'h02c9: q1 = 16'h2f00; // 0x0592
	13'h02ca: q1 = 16'h4eb9; // 0x0594
	13'h02cb: q1 = 16'h0000; // 0x0596
	13'h02cc: q1 = 16'h78f6; // 0x0598
	13'h02cd: q1 = 16'h4a9f; // 0x059a
	13'h02ce: q1 = 16'h200e; // 0x059c
	13'h02cf: q1 = 16'hd0bc; // 0x059e
	13'h02d0: q1 = 16'hffff; // 0x05a0
	13'h02d1: q1 = 16'hffe0; // 0x05a2
	13'h02d2: q1 = 16'h2e80; // 0x05a4
	13'h02d3: q1 = 16'h3f39; // 0x05a6
	13'h02d4: q1 = 16'h0001; // 0x05a8
	13'h02d5: q1 = 16'h8054; // 0x05aa
	13'h02d6: q1 = 16'h5257; // 0x05ac
	13'h02d7: q1 = 16'h4eb9; // 0x05ae
	13'h02d8: q1 = 16'h0000; // 0x05b0
	13'h02d9: q1 = 16'h0798; // 0x05b2
	13'h02da: q1 = 16'h4a5f; // 0x05b4
	13'h02db: q1 = 16'h0c79; // 0x05b6
	13'h02dc: q1 = 16'h0001; // 0x05b8
	13'h02dd: q1 = 16'h0001; // 0x05ba
	13'h02de: q1 = 16'h758c; // 0x05bc
	13'h02df: q1 = 16'h6618; // 0x05be
	13'h02e0: q1 = 16'h2ebc; // 0x05c0
	13'h02e1: q1 = 16'h0000; // 0x05c2
	13'h02e2: q1 = 16'hca10; // 0x05c4
	13'h02e3: q1 = 16'h200e; // 0x05c6
	13'h02e4: q1 = 16'hd0bc; // 0x05c8
	13'h02e5: q1 = 16'hffff; // 0x05ca
	13'h02e6: q1 = 16'hffe0; // 0x05cc
	13'h02e7: q1 = 16'h2f00; // 0x05ce
	13'h02e8: q1 = 16'h4eb9; // 0x05d0
	13'h02e9: q1 = 16'h0000; // 0x05d2
	13'h02ea: q1 = 16'h0770; // 0x05d4
	13'h02eb: q1 = 16'h4a9f; // 0x05d6
	13'h02ec: q1 = 16'h3e84; // 0x05d8
	13'h02ed: q1 = 16'h4267; // 0x05da
	13'h02ee: q1 = 16'h3f3c; // 0x05dc
	13'h02ef: q1 = 16'h0064; // 0x05de
	13'h02f0: q1 = 16'h3f3c; // 0x05e0
	13'h02f1: q1 = 16'h0011; // 0x05e2
	13'h02f2: q1 = 16'h200e; // 0x05e4
	13'h02f3: q1 = 16'hd0bc; // 0x05e6
	13'h02f4: q1 = 16'hffff; // 0x05e8
	13'h02f5: q1 = 16'hffe0; // 0x05ea
	13'h02f6: q1 = 16'h2f00; // 0x05ec
	13'h02f7: q1 = 16'h4eb9; // 0x05ee
	13'h02f8: q1 = 16'h0000; // 0x05f0
	13'h02f9: q1 = 16'h026c; // 0x05f2
	13'h02fa: q1 = 16'hdefc; // 0x05f4
	13'h02fb: q1 = 16'h000a; // 0x05f6
	13'h02fc: q1 = 16'hb87c; // 0x05f8
	13'h02fd: q1 = 16'h003f; // 0x05fa
	13'h02fe: q1 = 16'h6602; // 0x05fc
	13'h02ff: q1 = 16'h5245; // 0x05fe
	13'h0300: q1 = 16'hba7c; // 0x0600
	13'h0301: q1 = 16'h0003; // 0x0602
	13'h0302: q1 = 16'h671c; // 0x0604
	13'h0303: q1 = 16'h707d; // 0x0606
	13'h0304: q1 = 16'h9044; // 0x0608
	13'h0305: q1 = 16'h3800; // 0x060a
	13'h0306: q1 = 16'h33fc; // 0x060c
	13'h0307: q1 = 16'h0001; // 0x060e
	13'h0308: q1 = 16'h0001; // 0x0610
	13'h0309: q1 = 16'h86a8; // 0x0612
	13'h030a: q1 = 16'h4a79; // 0x0614
	13'h030b: q1 = 16'h0001; // 0x0616
	13'h030c: q1 = 16'h86a8; // 0x0618
	13'h030d: q1 = 16'h6702; // 0x061a
	13'h030e: q1 = 16'h60f6; // 0x061c
	13'h030f: q1 = 16'h6000; // 0x061e
	13'h0310: q1 = 16'hff66; // 0x0620
	13'h0311: q1 = 16'h3eb9; // 0x0622
	13'h0312: q1 = 16'h0001; // 0x0624
	13'h0313: q1 = 16'h8054; // 0x0626
	13'h0314: q1 = 16'h4eb9; // 0x0628
	13'h0315: q1 = 16'h0000; // 0x062a
	13'h0316: q1 = 16'ha9ae; // 0x062c
	13'h0317: q1 = 16'h2079; // 0x062e
	13'h0318: q1 = 16'h0001; // 0x0630
	13'h0319: q1 = 16'h7eb2; // 0x0632
	13'h031a: q1 = 16'h5250; // 0x0634
	13'h031b: q1 = 16'h2079; // 0x0636
	13'h031c: q1 = 16'h0001; // 0x0638
	13'h031d: q1 = 16'h7eb2; // 0x063a
	13'h031e: q1 = 16'h5368; // 0x063c
	13'h031f: q1 = 16'h0002; // 0x063e
	13'h0320: q1 = 16'h2079; // 0x0640
	13'h0321: q1 = 16'h0001; // 0x0642
	13'h0322: q1 = 16'h7eb2; // 0x0644
	13'h0323: q1 = 16'h5268; // 0x0646
	13'h0324: q1 = 16'h0004; // 0x0648
	13'h0325: q1 = 16'h2079; // 0x064a
	13'h0326: q1 = 16'h0001; // 0x064c
	13'h0327: q1 = 16'h7eb2; // 0x064e
	13'h0328: q1 = 16'h5368; // 0x0650
	13'h0329: q1 = 16'h0006; // 0x0652
	13'h032a: q1 = 16'h3c39; // 0x0654
	13'h032b: q1 = 16'h0001; // 0x0656
	13'h032c: q1 = 16'h862a; // 0x0658
	13'h032d: q1 = 16'h0c79; // 0x065a
	13'h032e: q1 = 16'h0002; // 0x065c
	13'h032f: q1 = 16'h0001; // 0x065e
	13'h0330: q1 = 16'h87dc; // 0x0660
	13'h0331: q1 = 16'h6606; // 0x0662
	13'h0332: q1 = 16'hdc79; // 0x0664
	13'h0333: q1 = 16'h0001; // 0x0666
	13'h0334: q1 = 16'h8650; // 0x0668
	13'h0335: q1 = 16'h4a46; // 0x066a
	13'h0336: q1 = 16'h6700; // 0x066c
	13'h0337: q1 = 16'h00c0; // 0x066e
	13'h0338: q1 = 16'h0c79; // 0x0670
	13'h0339: q1 = 16'h0001; // 0x0672
	13'h033a: q1 = 16'h0001; // 0x0674
	13'h033b: q1 = 16'h87dc; // 0x0676
	13'h033c: q1 = 16'h6700; // 0x0678
	13'h033d: q1 = 16'hfec2; // 0x067a
	13'h033e: q1 = 16'h3e39; // 0x067c
	13'h033f: q1 = 16'h0001; // 0x067e
	13'h0340: q1 = 16'h8054; // 0x0680
	13'h0341: q1 = 16'h7001; // 0x0682
	13'h0342: q1 = 16'h9079; // 0x0684
	13'h0343: q1 = 16'h0001; // 0x0686
	13'h0344: q1 = 16'h8054; // 0x0688
	13'h0345: q1 = 16'h33c0; // 0x068a
	13'h0346: q1 = 16'h0001; // 0x068c
	13'h0347: q1 = 16'h8054; // 0x068e
	13'h0348: q1 = 16'h3039; // 0x0690
	13'h0349: q1 = 16'h0001; // 0x0692
	13'h034a: q1 = 16'h8054; // 0x0694
	13'h034b: q1 = 16'hc1fc; // 0x0696
	13'h034c: q1 = 16'h0026; // 0x0698
	13'h034d: q1 = 16'hd0bc; // 0x069a
	13'h034e: q1 = 16'h0001; // 0x069c
	13'h034f: q1 = 16'h862a; // 0x069e
	13'h0350: q1 = 16'h2040; // 0x06a0
	13'h0351: q1 = 16'h4a50; // 0x06a2
	13'h0352: q1 = 16'h660e; // 0x06a4
	13'h0353: q1 = 16'h7001; // 0x06a6
	13'h0354: q1 = 16'h9079; // 0x06a8
	13'h0355: q1 = 16'h0001; // 0x06aa
	13'h0356: q1 = 16'h8054; // 0x06ac
	13'h0357: q1 = 16'h33c0; // 0x06ae
	13'h0358: q1 = 16'h0001; // 0x06b0
	13'h0359: q1 = 16'h8054; // 0x06b2
	13'h035a: q1 = 16'h3039; // 0x06b4
	13'h035b: q1 = 16'h0001; // 0x06b6
	13'h035c: q1 = 16'h8054; // 0x06b8
	13'h035d: q1 = 16'hc1fc; // 0x06ba
	13'h035e: q1 = 16'h0026; // 0x06bc
	13'h035f: q1 = 16'hd0bc; // 0x06be
	13'h0360: q1 = 16'h0001; // 0x06c0
	13'h0361: q1 = 16'h8628; // 0x06c2
	13'h0362: q1 = 16'h23c0; // 0x06c4
	13'h0363: q1 = 16'h0001; // 0x06c6
	13'h0364: q1 = 16'h7fb8; // 0x06c8
	13'h0365: q1 = 16'h4eb9; // 0x06ca
	13'h0366: q1 = 16'h0000; // 0x06cc
	13'h0367: q1 = 16'h0226; // 0x06ce
	13'h0368: q1 = 16'h0c79; // 0x06d0
	13'h0369: q1 = 16'h0001; // 0x06d2
	13'h036a: q1 = 16'h0001; // 0x06d4
	13'h036b: q1 = 16'h8054; // 0x06d6
	13'h036c: q1 = 16'h6618; // 0x06d8
	13'h036d: q1 = 16'h4a79; // 0x06da
	13'h036e: q1 = 16'h0001; // 0x06dc
	13'h036f: q1 = 16'h758e; // 0x06de
	13'h0370: q1 = 16'h6710; // 0x06e0
	13'h0371: q1 = 16'h33fc; // 0x06e2
	13'h0372: q1 = 16'h0001; // 0x06e4
	13'h0373: q1 = 16'h0001; // 0x06e6
	13'h0374: q1 = 16'h7fa6; // 0x06e8
	13'h0375: q1 = 16'h33fc; // 0x06ea
	13'h0376: q1 = 16'h0001; // 0x06ec
	13'h0377: q1 = 16'h0001; // 0x06ee
	13'h0378: q1 = 16'h8052; // 0x06f0
	13'h0379: q1 = 16'h4a79; // 0x06f2
	13'h037a: q1 = 16'h0001; // 0x06f4
	13'h037b: q1 = 16'h8054; // 0x06f6
	13'h037c: q1 = 16'h6614; // 0x06f8
	13'h037d: q1 = 16'h4a79; // 0x06fa
	13'h037e: q1 = 16'h0001; // 0x06fc
	13'h037f: q1 = 16'h758e; // 0x06fe
	13'h0380: q1 = 16'h670c; // 0x0700
	13'h0381: q1 = 16'h4279; // 0x0702
	13'h0382: q1 = 16'h0001; // 0x0704
	13'h0383: q1 = 16'h7fa6; // 0x0706
	13'h0384: q1 = 16'h4279; // 0x0708
	13'h0385: q1 = 16'h0001; // 0x070a
	13'h0386: q1 = 16'h8052; // 0x070c
	13'h0387: q1 = 16'hbe79; // 0x070e
	13'h0388: q1 = 16'h0001; // 0x0710
	13'h0389: q1 = 16'h8054; // 0x0712
	13'h038a: q1 = 16'h6714; // 0x0714
	13'h038b: q1 = 16'h33fc; // 0x0716
	13'h038c: q1 = 16'h0001; // 0x0718
	13'h038d: q1 = 16'h0001; // 0x071a
	13'h038e: q1 = 16'h7fc8; // 0x071c
	13'h038f: q1 = 16'h3eb9; // 0x071e
	13'h0390: q1 = 16'h0001; // 0x0720
	13'h0391: q1 = 16'h8054; // 0x0722
	13'h0392: q1 = 16'h4eb9; // 0x0724
	13'h0393: q1 = 16'h0000; // 0x0726
	13'h0394: q1 = 16'had5a; // 0x0728
	13'h0395: q1 = 16'h6000; // 0x072a
	13'h0396: q1 = 16'hfe10; // 0x072c
	13'h0397: q1 = 16'h4a9f; // 0x072e
	13'h0398: q1 = 16'h4cdf; // 0x0730
	13'h0399: q1 = 16'h00f0; // 0x0732
	13'h039a: q1 = 16'h4e5e; // 0x0734
	13'h039b: q1 = 16'h4e75; // 0x0736
	13'h039c: q1 = 16'h4e56; // 0x0738
	13'h039d: q1 = 16'h0000; // 0x073a
	13'h039e: q1 = 16'h48e7; // 0x073c
	13'h039f: q1 = 16'h0104; // 0x073e
	13'h03a0: q1 = 16'h2a7c; // 0x0740
	13'h03a1: q1 = 16'h0001; // 0x0742
	13'h03a2: q1 = 16'h7f2c; // 0x0744
	13'h03a3: q1 = 16'h302d; // 0x0746
	13'h03a4: q1 = 16'h0018; // 0x0748
	13'h03a5: q1 = 16'h4a9f; // 0x074a
	13'h03a6: q1 = 16'h4cdf; // 0x074c
	13'h03a7: q1 = 16'h2000; // 0x074e
	13'h03a8: q1 = 16'h4e5e; // 0x0750
	13'h03a9: q1 = 16'h4e75; // 0x0752
	13'h03aa: q1 = 16'h4e56; // 0x0754
	13'h03ab: q1 = 16'h0000; // 0x0756
	13'h03ac: q1 = 16'h48e7; // 0x0758
	13'h03ad: q1 = 16'h0104; // 0x075a
	13'h03ae: q1 = 16'h2a7c; // 0x075c
	13'h03af: q1 = 16'h0001; // 0x075e
	13'h03b0: q1 = 16'h7f2c; // 0x0760
	13'h03b1: q1 = 16'h42ad; // 0x0762
	13'h03b2: q1 = 16'h0006; // 0x0764
	13'h03b3: q1 = 16'h4a9f; // 0x0766
	13'h03b4: q1 = 16'h4cdf; // 0x0768
	13'h03b5: q1 = 16'h2000; // 0x076a
	13'h03b6: q1 = 16'h4e5e; // 0x076c
	13'h03b7: q1 = 16'h4e75; // 0x076e
	13'h03b8: q1 = 16'h4e56; // 0x0770
	13'h03b9: q1 = 16'h0000; // 0x0772
	13'h03ba: q1 = 16'h48e7; // 0x0774
	13'h03bb: q1 = 16'h0104; // 0x0776
	13'h03bc: q1 = 16'h2a7c; // 0x0778
	13'h03bd: q1 = 16'h0001; // 0x077a
	13'h03be: q1 = 16'h7f2c; // 0x077c
	13'h03bf: q1 = 16'h4a6e; // 0x077e
	13'h03c0: q1 = 16'h0008; // 0x0780
	13'h03c1: q1 = 16'h662e; // 0x0782
	13'h03c2: q1 = 16'h3b7c; // 0x0784
	13'h03c3: q1 = 16'h0001; // 0x0786
	13'h03c4: q1 = 16'h001a; // 0x0788
	13'h03c5: q1 = 16'h3b7c; // 0x078a
	13'h03c6: q1 = 16'h0001; // 0x078c
	13'h03c7: q1 = 16'h0018; // 0x078e
	13'h03c8: q1 = 16'h23fc; // 0x0790
	13'h03c9: q1 = 16'h0000; // 0x0792
	13'h03ca: q1 = 16'hccb0; // 0x0794
	13'h03cb: q1 = 16'h0001; // 0x0796
	13'h03cc: q1 = 16'h86ae; // 0x0798
	13'h03cd: q1 = 16'h23fc; // 0x079a
	13'h03ce: q1 = 16'h0000; // 0x079c
	13'h03cf: q1 = 16'hce3a; // 0x079e
	13'h03d0: q1 = 16'h0001; // 0x07a0
	13'h03d1: q1 = 16'h7ebc; // 0x07a2
	13'h03d2: q1 = 16'h4279; // 0x07a4
	13'h03d3: q1 = 16'h0001; // 0x07a6
	13'h03d4: q1 = 16'h7ba2; // 0x07a8
	13'h03d5: q1 = 16'h4279; // 0x07aa
	13'h03d6: q1 = 16'h0001; // 0x07ac
	13'h03d7: q1 = 16'h7ba4; // 0x07ae
	13'h03d8: q1 = 16'h602c; // 0x07b0
	13'h03d9: q1 = 16'h0c6e; // 0x07b2
	13'h03da: q1 = 16'h0001; // 0x07b4
	13'h03db: q1 = 16'h0008; // 0x07b6
	13'h03dc: q1 = 16'h6624; // 0x07b8
	13'h03dd: q1 = 16'h206d; // 0x07ba
	13'h03de: q1 = 16'h0024; // 0x07bc
	13'h03df: q1 = 16'h30bc; // 0x07be
	13'h03e0: q1 = 16'h0080; // 0x07c0
	13'h03e1: q1 = 16'h206d; // 0x07c2
	13'h03e2: q1 = 16'h0024; // 0x07c4
	13'h03e3: q1 = 16'h317c; // 0x07c6
	13'h03e4: q1 = 16'h1800; // 0x07c8
	13'h03e5: q1 = 16'h0002; // 0x07ca
	13'h03e6: q1 = 16'h426d; // 0x07cc
	13'h03e7: q1 = 16'h000e; // 0x07ce
	13'h03e8: q1 = 16'h42ad; // 0x07d0
	13'h03e9: q1 = 16'h0006; // 0x07d2
	13'h03ea: q1 = 16'h4eb9; // 0x07d4
	13'h03eb: q1 = 16'h0000; // 0x07d6
	13'h03ec: q1 = 16'h61f8; // 0x07d8
	13'h03ed: q1 = 16'h3abc; // 0x07da
	13'h03ee: q1 = 16'h0001; // 0x07dc
	13'h03ef: q1 = 16'h4a9f; // 0x07de
	13'h03f0: q1 = 16'h4cdf; // 0x07e0
	13'h03f1: q1 = 16'h2000; // 0x07e2
	13'h03f2: q1 = 16'h4e5e; // 0x07e4
	13'h03f3: q1 = 16'h4e75; // 0x07e6
	13'h03f4: q1 = 16'h4e56; // 0x07e8
	13'h03f5: q1 = 16'h0000; // 0x07ea
	13'h03f6: q1 = 16'h48e7; // 0x07ec
	13'h03f7: q1 = 16'h0104; // 0x07ee
	13'h03f8: q1 = 16'h2a7c; // 0x07f0
	13'h03f9: q1 = 16'h0001; // 0x07f2
	13'h03fa: q1 = 16'h7f2c; // 0x07f4
	13'h03fb: q1 = 16'h206d; // 0x07f6
	13'h03fc: q1 = 16'h0024; // 0x07f8
	13'h03fd: q1 = 16'h30bc; // 0x07fa
	13'h03fe: q1 = 16'h3c00; // 0x07fc
	13'h03ff: q1 = 16'h206d; // 0x07fe
	13'h0400: q1 = 16'h0024; // 0x0800
	13'h0401: q1 = 16'h317c; // 0x0802
	13'h0402: q1 = 16'h4080; // 0x0804
	13'h0403: q1 = 16'h0002; // 0x0806
	13'h0404: q1 = 16'h426d; // 0x0808
	13'h0405: q1 = 16'h000e; // 0x080a
	13'h0406: q1 = 16'h42ad; // 0x080c
	13'h0407: q1 = 16'h0006; // 0x080e
	13'h0408: q1 = 16'h4eb9; // 0x0810
	13'h0409: q1 = 16'h0000; // 0x0812
	13'h040a: q1 = 16'h61f8; // 0x0814
	13'h040b: q1 = 16'h4a9f; // 0x0816
	13'h040c: q1 = 16'h4cdf; // 0x0818
	13'h040d: q1 = 16'h2000; // 0x081a
	13'h040e: q1 = 16'h4e5e; // 0x081c
	13'h040f: q1 = 16'h4e75; // 0x081e
	13'h0410: q1 = 16'h4e56; // 0x0820
	13'h0411: q1 = 16'hfff4; // 0x0822
	13'h0412: q1 = 16'h48e7; // 0x0824
	13'h0413: q1 = 16'h3f1c; // 0x0826
	13'h0414: q1 = 16'h2a7c; // 0x0828
	13'h0415: q1 = 16'h0001; // 0x082a
	13'h0416: q1 = 16'h7f2c; // 0x082c
	13'h0417: q1 = 16'h4aad; // 0x082e
	13'h0418: q1 = 16'h001c; // 0x0830
	13'h0419: q1 = 16'h6f04; // 0x0832
	13'h041a: q1 = 16'h53ad; // 0x0834
	13'h041b: q1 = 16'h001c; // 0x0836
	13'h041c: q1 = 16'h4a6d; // 0x0838
	13'h041d: q1 = 16'h0018; // 0x083a
	13'h041e: q1 = 16'h6600; // 0x083c
	13'h041f: q1 = 16'h0536; // 0x083e
	13'h0420: q1 = 16'h4a6d; // 0x0840
	13'h0421: q1 = 16'h001a; // 0x0842
	13'h0422: q1 = 16'h6720; // 0x0844
	13'h0423: q1 = 16'h0c6d; // 0x0846
	13'h0424: q1 = 16'h0005; // 0x0848
	13'h0425: q1 = 16'h001a; // 0x084a
	13'h0426: q1 = 16'h6718; // 0x084c
	13'h0427: q1 = 16'h4eb9; // 0x084e
	13'h0428: q1 = 16'h0000; // 0x0850
	13'h0429: q1 = 16'h524a; // 0x0852
	13'h042a: q1 = 16'h0c6d; // 0x0854
	13'h042b: q1 = 16'h0004; // 0x0856
	13'h042c: q1 = 16'h001a; // 0x0858
	13'h042d: q1 = 16'h6600; // 0x085a
	13'h042e: q1 = 16'h04c8; // 0x085c
	13'h042f: q1 = 16'h4a6d; // 0x085e
	13'h0430: q1 = 16'h0018; // 0x0860
	13'h0431: q1 = 16'h6600; // 0x0862
	13'h0432: q1 = 16'h04c0; // 0x0864
	13'h0433: q1 = 16'h0c6d; // 0x0866
	13'h0434: q1 = 16'h0005; // 0x0868
	13'h0435: q1 = 16'h001a; // 0x086a
	13'h0436: q1 = 16'h6622; // 0x086c
	13'h0437: q1 = 16'h4a79; // 0x086e
	13'h0438: q1 = 16'h0001; // 0x0870
	13'h0439: q1 = 16'h7fc6; // 0x0872
	13'h043a: q1 = 16'h6704; // 0x0874
	13'h043b: q1 = 16'h7e01; // 0x0876
	13'h043c: q1 = 16'h6008; // 0x0878
	13'h043d: q1 = 16'h4eb9; // 0x087a
	13'h043e: q1 = 16'h0000; // 0x087c
	13'h043f: q1 = 16'h5688; // 0x087e
	13'h0440: q1 = 16'h3e00; // 0x0880
	13'h0441: q1 = 16'h4a47; // 0x0882
	13'h0442: q1 = 16'h6706; // 0x0884
	13'h0443: q1 = 16'h3b7c; // 0x0886
	13'h0444: q1 = 16'h0002; // 0x0888
	13'h0445: q1 = 16'h0018; // 0x088a
	13'h0446: q1 = 16'h6000; // 0x088c
	13'h0447: q1 = 16'h04e6; // 0x088e
	13'h0448: q1 = 16'h4257; // 0x0890
	13'h0449: q1 = 16'h206d; // 0x0892
	13'h044a: q1 = 16'h0024; // 0x0894
	13'h044b: q1 = 16'h3f28; // 0x0896
	13'h044c: q1 = 16'h0002; // 0x0898
	13'h044d: q1 = 16'h206d; // 0x089a
	13'h044e: q1 = 16'h0024; // 0x089c
	13'h044f: q1 = 16'h3f10; // 0x089e
	13'h0450: q1 = 16'h4eb9; // 0x08a0
	13'h0451: q1 = 16'h0000; // 0x08a2
	13'h0452: q1 = 16'h42d4; // 0x08a4
	13'h0453: q1 = 16'h4a9f; // 0x08a6
	13'h0454: q1 = 16'h4a40; // 0x08a8
	13'h0455: q1 = 16'h671a; // 0x08aa
	13'h0456: q1 = 16'h0c6d; // 0x08ac
	13'h0457: q1 = 16'h0004; // 0x08ae
	13'h0458: q1 = 16'h001a; // 0x08b0
	13'h0459: q1 = 16'h6712; // 0x08b2
	13'h045a: q1 = 16'h4255; // 0x08b4
	13'h045b: q1 = 16'h3b7c; // 0x08b6
	13'h045c: q1 = 16'h0024; // 0x08b8
	13'h045d: q1 = 16'h000e; // 0x08ba
	13'h045e: q1 = 16'h3b7c; // 0x08bc
	13'h045f: q1 = 16'h0005; // 0x08be
	13'h0460: q1 = 16'h001a; // 0x08c0
	13'h0461: q1 = 16'h6000; // 0x08c2
	13'h0462: q1 = 16'h04b0; // 0x08c4
	13'h0463: q1 = 16'h0c6d; // 0x08c6
	13'h0464: q1 = 16'h0004; // 0x08c8
	13'h0465: q1 = 16'h001a; // 0x08ca
	13'h0466: q1 = 16'h6714; // 0x08cc
	13'h0467: q1 = 16'h4a79; // 0x08ce
	13'h0468: q1 = 16'h0001; // 0x08d0
	13'h0469: q1 = 16'h7f20; // 0x08d2
	13'h046a: q1 = 16'h660c; // 0x08d4
	13'h046b: q1 = 16'h4eb9; // 0x08d6
	13'h046c: q1 = 16'h0000; // 0x08d8
	13'h046d: q1 = 16'h4f80; // 0x08da
	13'h046e: q1 = 16'h4a40; // 0x08dc
	13'h046f: q1 = 16'h6600; // 0x08de
	13'h0470: q1 = 16'h0444; // 0x08e0
	13'h0471: q1 = 16'h3839; // 0x08e2
	13'h0472: q1 = 16'h0001; // 0x08e4
	13'h0473: q1 = 16'h8622; // 0x08e6
	13'h0474: q1 = 16'h3639; // 0x08e8
	13'h0475: q1 = 16'h0001; // 0x08ea
	13'h0476: q1 = 16'h8624; // 0x08ec
	13'h0477: q1 = 16'h4a79; // 0x08ee
	13'h0478: q1 = 16'h0001; // 0x08f0
	13'h0479: q1 = 16'h7fc6; // 0x08f2
	13'h047a: q1 = 16'h6712; // 0x08f4
	13'h047b: q1 = 16'h4a79; // 0x08f6
	13'h047c: q1 = 16'h0001; // 0x08f8
	13'h047d: q1 = 16'h806e; // 0x08fa
	13'h047e: q1 = 16'h660a; // 0x08fc
	13'h047f: q1 = 16'h3b79; // 0x08fe
	13'h0480: q1 = 16'h0001; // 0x0900
	13'h0481: q1 = 16'h8682; // 0x0902
	13'h0482: q1 = 16'h000e; // 0x0904
	13'h0483: q1 = 16'h6030; // 0x0906
	13'h0484: q1 = 16'h4a79; // 0x0908
	13'h0485: q1 = 16'h0001; // 0x090a
	13'h0486: q1 = 16'h7b9e; // 0x090c
	13'h0487: q1 = 16'h6710; // 0x090e
	13'h0488: q1 = 16'h4a79; // 0x0910
	13'h0489: q1 = 16'h0001; // 0x0912
	13'h048a: q1 = 16'h8676; // 0x0914
	13'h048b: q1 = 16'h6708; // 0x0916
	13'h048c: q1 = 16'h3b7c; // 0x0918
	13'h048d: q1 = 16'h0024; // 0x091a
	13'h048e: q1 = 16'h000e; // 0x091c
	13'h048f: q1 = 16'h6018; // 0x091e
	13'h0490: q1 = 16'h0c6d; // 0x0920
	13'h0491: q1 = 16'h0004; // 0x0922
	13'h0492: q1 = 16'h001a; // 0x0924
	13'h0493: q1 = 16'h6710; // 0x0926
	13'h0494: q1 = 16'h3e83; // 0x0928
	13'h0495: q1 = 16'h3f04; // 0x092a
	13'h0496: q1 = 16'h4eb9; // 0x092c
	13'h0497: q1 = 16'h0000; // 0x092e
	13'h0498: q1 = 16'h0a1c; // 0x0930
	13'h0499: q1 = 16'h4a5f; // 0x0932
	13'h049a: q1 = 16'h3b40; // 0x0934
	13'h049b: q1 = 16'h000e; // 0x0936
	13'h049c: q1 = 16'h4a79; // 0x0938
	13'h049d: q1 = 16'h0001; // 0x093a
	13'h049e: q1 = 16'h7fc6; // 0x093c
	13'h049f: q1 = 16'h6714; // 0x093e
	13'h04a0: q1 = 16'h4a79; // 0x0940
	13'h04a1: q1 = 16'h0001; // 0x0942
	13'h04a2: q1 = 16'h806e; // 0x0944
	13'h04a3: q1 = 16'h660c; // 0x0946
	13'h04a4: q1 = 16'h3d79; // 0x0948
	13'h04a5: q1 = 16'h0001; // 0x094a
	13'h04a6: q1 = 16'h8880; // 0x094c
	13'h04a7: q1 = 16'hfffa; // 0x094e
	13'h04a8: q1 = 16'h6000; // 0x0950
	13'h04a9: q1 = 16'h0096; // 0x0952
	13'h04aa: q1 = 16'h0c6d; // 0x0954
	13'h04ab: q1 = 16'h0004; // 0x0956
	13'h04ac: q1 = 16'h001a; // 0x0958
	13'h04ad: q1 = 16'h660a; // 0x095a
	13'h04ae: q1 = 16'h3d7c; // 0x095c
	13'h04af: q1 = 16'h0001; // 0x095e
	13'h04b0: q1 = 16'hfffa; // 0x0960
	13'h04b1: q1 = 16'h6000; // 0x0962
	13'h04b2: q1 = 16'h0084; // 0x0964
	13'h04b3: q1 = 16'h4a79; // 0x0966
	13'h04b4: q1 = 16'h0001; // 0x0968
	13'h04b5: q1 = 16'h7b9e; // 0x096a
	13'h04b6: q1 = 16'h6608; // 0x096c
	13'h04b7: q1 = 16'h4a79; // 0x096e
	13'h04b8: q1 = 16'h0001; // 0x0970
	13'h04b9: q1 = 16'h7f20; // 0x0972
	13'h04ba: q1 = 16'h6706; // 0x0974
	13'h04bb: q1 = 16'h426e; // 0x0976
	13'h04bc: q1 = 16'hfffa; // 0x0978
	13'h04bd: q1 = 16'h606c; // 0x097a
	13'h04be: q1 = 16'h2079; // 0x097c
	13'h04bf: q1 = 16'h0001; // 0x097e
	13'h04c0: q1 = 16'h7eb2; // 0x0980
	13'h04c1: q1 = 16'h3f28; // 0x0982
	13'h04c2: q1 = 16'h0006; // 0x0984
	13'h04c3: q1 = 16'h2079; // 0x0986
	13'h04c4: q1 = 16'h0001; // 0x0988
	13'h04c5: q1 = 16'h7eb2; // 0x098a
	13'h04c6: q1 = 16'h3028; // 0x098c
	13'h04c7: q1 = 16'h0004; // 0x098e
	13'h04c8: q1 = 16'h9157; // 0x0990
	13'h04c9: q1 = 16'h2079; // 0x0992
	13'h04ca: q1 = 16'h0001; // 0x0994
	13'h04cb: q1 = 16'h7eb2; // 0x0996
	13'h04cc: q1 = 16'h3028; // 0x0998
	13'h04cd: q1 = 16'h0002; // 0x099a
	13'h04ce: q1 = 16'h2279; // 0x099c
	13'h04cf: q1 = 16'h0001; // 0x099e
	13'h04d0: q1 = 16'h7eb2; // 0x09a0
	13'h04d1: q1 = 16'h9051; // 0x09a2
	13'h04d2: q1 = 16'hd05f; // 0x09a4
	13'h04d3: q1 = 16'h3e00; // 0x09a6
	13'h04d4: q1 = 16'he247; // 0x09a8
	13'h04d5: q1 = 16'h3007; // 0x09aa
	13'h04d6: q1 = 16'he240; // 0x09ac
	13'h04d7: q1 = 16'h3207; // 0x09ae
	13'h04d8: q1 = 16'he641; // 0x09b0
	13'h04d9: q1 = 16'h9041; // 0x09b2
	13'h04da: q1 = 16'h3a00; // 0x09b4
	13'h04db: q1 = 16'h4a44; // 0x09b6
	13'h04dc: q1 = 16'h6c06; // 0x09b8
	13'h04dd: q1 = 16'h3004; // 0x09ba
	13'h04de: q1 = 16'h4440; // 0x09bc
	13'h04df: q1 = 16'h3800; // 0x09be
	13'h04e0: q1 = 16'h4a43; // 0x09c0
	13'h04e1: q1 = 16'h6c06; // 0x09c2
	13'h04e2: q1 = 16'h3003; // 0x09c4
	13'h04e3: q1 = 16'h4440; // 0x09c6
	13'h04e4: q1 = 16'h3600; // 0x09c8
	13'h04e5: q1 = 16'hb843; // 0x09ca
	13'h04e6: q1 = 16'h6f04; // 0x09cc
	13'h04e7: q1 = 16'he243; // 0x09ce
	13'h04e8: q1 = 16'h6002; // 0x09d0
	13'h04e9: q1 = 16'he244; // 0x09d2
	13'h04ea: q1 = 16'h3004; // 0x09d4
	13'h04eb: q1 = 16'hd043; // 0x09d6
	13'h04ec: q1 = 16'hb045; // 0x09d8
	13'h04ed: q1 = 16'h6f08; // 0x09da
	13'h04ee: q1 = 16'h3d7c; // 0x09dc
	13'h04ef: q1 = 16'h0001; // 0x09de
	13'h04f0: q1 = 16'hfffa; // 0x09e0
	13'h04f1: q1 = 16'h6004; // 0x09e2
	13'h04f2: q1 = 16'h426e; // 0x09e4
	13'h04f3: q1 = 16'hfffa; // 0x09e6
	13'h04f4: q1 = 16'h4a79; // 0x09e8
	13'h04f5: q1 = 16'h0001; // 0x09ea
	13'h04f6: q1 = 16'h7fc6; // 0x09ec
	13'h04f7: q1 = 16'h6712; // 0x09ee
	13'h04f8: q1 = 16'h4a79; // 0x09f0
	13'h04f9: q1 = 16'h0001; // 0x09f2
	13'h04fa: q1 = 16'h806e; // 0x09f4
	13'h04fb: q1 = 16'h660a; // 0x09f6
	13'h04fc: q1 = 16'h3d79; // 0x09f8
	13'h04fd: q1 = 16'h0001; // 0x09fa
	13'h04fe: q1 = 16'h81fa; // 0x09fc
	13'h04ff: q1 = 16'hfff8; // 0x09fe
	13'h0500: q1 = 16'h6026; // 0x0a00
	13'h0501: q1 = 16'h4a79; // 0x0a02
	13'h0502: q1 = 16'h0001; // 0x0a04
	13'h0503: q1 = 16'h7b9e; // 0x0a06
	13'h0504: q1 = 16'h6706; // 0x0a08
	13'h0505: q1 = 16'h426e; // 0x0a0a
	13'h0506: q1 = 16'hfff8; // 0x0a0c
	13'h0507: q1 = 16'h6018; // 0x0a0e
	13'h0508: q1 = 16'h4a79; // 0x0a10
	13'h0509: q1 = 16'h0001; // 0x0a12
	13'h050a: q1 = 16'h7f20; // 0x0a14
	13'h050b: q1 = 16'h6708; // 0x0a16
	13'h050c: q1 = 16'h3d7c; // 0x0a18
	13'h050d: q1 = 16'h0001; // 0x0a1a
	13'h050e: q1 = 16'hfff8; // 0x0a1c
	13'h050f: q1 = 16'h6008; // 0x0a1e
	13'h0510: q1 = 16'h3d79; // 0x0a20
	13'h0511: q1 = 16'h0001; // 0x0a22
	13'h0512: q1 = 16'h7fca; // 0x0a24
	13'h0513: q1 = 16'hfff8; // 0x0a26
	13'h0514: q1 = 16'h4a79; // 0x0a28
	13'h0515: q1 = 16'h0001; // 0x0a2a
	13'h0516: q1 = 16'h7590; // 0x0a2c
	13'h0517: q1 = 16'h673e; // 0x0a2e
	13'h0518: q1 = 16'h42ae; // 0x0a30
	13'h0519: q1 = 16'hfff4; // 0x0a32
	13'h051a: q1 = 16'h2039; // 0x0a34
	13'h051b: q1 = 16'h0000; // 0x0a36
	13'h051c: q1 = 16'hcafe; // 0x0a38
	13'h051d: q1 = 16'he580; // 0x0a3a
	13'h051e: q1 = 16'hd1ae; // 0x0a3c
	13'h051f: q1 = 16'hfff4; // 0x0a3e
	13'h0520: q1 = 16'h202e; // 0x0a40
	13'h0521: q1 = 16'hfff4; // 0x0a42
	13'h0522: q1 = 16'he680; // 0x0a44
	13'h0523: q1 = 16'h2d40; // 0x0a46
	13'h0524: q1 = 16'hfff4; // 0x0a48
	13'h0525: q1 = 16'h206e; // 0x0a4a
	13'h0526: q1 = 16'hfff4; // 0x0a4c
	13'h0527: q1 = 16'h2010; // 0x0a4e
	13'h0528: q1 = 16'he880; // 0x0a50
	13'h0529: q1 = 16'hb0b9; // 0x0a52
	13'h052a: q1 = 16'h0000; // 0x0a54
	13'h052b: q1 = 16'hcb02; // 0x0a56
	13'h052c: q1 = 16'h6614; // 0x0a58
	13'h052d: q1 = 16'h206e; // 0x0a5a
	13'h052e: q1 = 16'hfff4; // 0x0a5c
	13'h052f: q1 = 16'h317c; // 0x0a5e
	13'h0530: q1 = 16'h000a; // 0x0a60
	13'h0531: q1 = 16'hffe4; // 0x0a62
	13'h0532: q1 = 16'h7014; // 0x0a64
	13'h0533: q1 = 16'h226e; // 0x0a66
	13'h0534: q1 = 16'hfff4; // 0x0a68
	13'h0535: q1 = 16'hd169; // 0x0a6a
	13'h0536: q1 = 16'hffe4; // 0x0a6c
	13'h0537: q1 = 16'h4a79; // 0x0a6e
	13'h0538: q1 = 16'h0001; // 0x0a70
	13'h0539: q1 = 16'h7fc6; // 0x0a72
	13'h053a: q1 = 16'h6708; // 0x0a74
	13'h053b: q1 = 16'h4a79; // 0x0a76
	13'h053c: q1 = 16'h0001; // 0x0a78
	13'h053d: q1 = 16'h806e; // 0x0a7a
	13'h053e: q1 = 16'h673e; // 0x0a7c
	13'h053f: q1 = 16'h4a79; // 0x0a7e
	13'h0540: q1 = 16'h0001; // 0x0a80
	13'h0541: q1 = 16'h7b9e; // 0x0a82
	13'h0542: q1 = 16'h6636; // 0x0a84
	13'h0543: q1 = 16'h4a79; // 0x0a86
	13'h0544: q1 = 16'h0001; // 0x0a88
	13'h0545: q1 = 16'h7f20; // 0x0a8a
	13'h0546: q1 = 16'h662e; // 0x0a8c
	13'h0547: q1 = 16'h0c6d; // 0x0a8e
	13'h0548: q1 = 16'h0004; // 0x0a90
	13'h0549: q1 = 16'h001a; // 0x0a92
	13'h054a: q1 = 16'h6726; // 0x0a94
	13'h054b: q1 = 16'h200e; // 0x0a96
	13'h054c: q1 = 16'hd0bc; // 0x0a98
	13'h054d: q1 = 16'hffff; // 0x0a9a
	13'h054e: q1 = 16'hfffa; // 0x0a9c
	13'h054f: q1 = 16'h2e80; // 0x0a9e
	13'h0550: q1 = 16'h200e; // 0x0aa0
	13'h0551: q1 = 16'hd0bc; // 0x0aa2
	13'h0552: q1 = 16'hffff; // 0x0aa4
	13'h0553: q1 = 16'hfff8; // 0x0aa6
	13'h0554: q1 = 16'h2f00; // 0x0aa8
	13'h0555: q1 = 16'h200d; // 0x0aaa
	13'h0556: q1 = 16'hd0bc; // 0x0aac
	13'h0557: q1 = 16'h0000; // 0x0aae
	13'h0558: q1 = 16'h000e; // 0x0ab0
	13'h0559: q1 = 16'h2f00; // 0x0ab2
	13'h055a: q1 = 16'h4eb9; // 0x0ab4
	13'h055b: q1 = 16'h0000; // 0x0ab6
	13'h055c: q1 = 16'h5f56; // 0x0ab8
	13'h055d: q1 = 16'hbf8f; // 0x0aba
	13'h055e: q1 = 16'h4a6e; // 0x0abc
	13'h055f: q1 = 16'hfffa; // 0x0abe
	13'h0560: q1 = 16'h6606; // 0x0ac0
	13'h0561: q1 = 16'h426d; // 0x0ac2
	13'h0562: q1 = 16'h0010; // 0x0ac4
	13'h0563: q1 = 16'h6034; // 0x0ac6
	13'h0564: q1 = 16'h0c6d; // 0x0ac8
	13'h0565: q1 = 16'h0004; // 0x0aca
	13'h0566: q1 = 16'h001a; // 0x0acc
	13'h0567: q1 = 16'h672c; // 0x0ace
	13'h0568: q1 = 16'h2079; // 0x0ad0
	13'h0569: q1 = 16'h0001; // 0x0ad2
	13'h056a: q1 = 16'h7fb8; // 0x0ad4
	13'h056b: q1 = 16'h3010; // 0x0ad6
	13'h056c: q1 = 16'h5340; // 0x0ad8
	13'h056d: q1 = 16'he740; // 0x0ada
	13'h056e: q1 = 16'hd07c; // 0x0adc
	13'h056f: q1 = 16'h00bc; // 0x0ade
	13'h0570: q1 = 16'h3b40; // 0x0ae0
	13'h0571: q1 = 16'h0010; // 0x0ae2
	13'h0572: q1 = 16'h2079; // 0x0ae4
	13'h0573: q1 = 16'h0001; // 0x0ae6
	13'h0574: q1 = 16'h7fb8; // 0x0ae8
	13'h0575: q1 = 16'h0c50; // 0x0aea
	13'h0576: q1 = 16'h0032; // 0x0aec
	13'h0577: q1 = 16'h6c08; // 0x0aee
	13'h0578: q1 = 16'h3b7c; // 0x0af0
	13'h0579: q1 = 16'h0001; // 0x0af2
	13'h057a: q1 = 16'h0004; // 0x0af4
	13'h057b: q1 = 16'h6004; // 0x0af6
	13'h057c: q1 = 16'h426d; // 0x0af8
	13'h057d: q1 = 16'h0004; // 0x0afa
	13'h057e: q1 = 16'h4a6d; // 0x0afc
	13'h057f: q1 = 16'h0010; // 0x0afe
	13'h0580: q1 = 16'h6700; // 0x0b00
	13'h0581: q1 = 16'h0122; // 0x0b02
	13'h0582: q1 = 16'h426e; // 0x0b04
	13'h0583: q1 = 16'hfffe; // 0x0b06
	13'h0584: q1 = 16'h426e; // 0x0b08
	13'h0585: q1 = 16'hfffc; // 0x0b0a
	13'h0586: q1 = 16'h3ead; // 0x0b0c
	13'h0587: q1 = 16'h0010; // 0x0b0e
	13'h0588: q1 = 16'h3f2d; // 0x0b10
	13'h0589: q1 = 16'h000e; // 0x0b12
	13'h058a: q1 = 16'h4eb9; // 0x0b14
	13'h058b: q1 = 16'h0000; // 0x0b16
	13'h058c: q1 = 16'h1280; // 0x0b18
	13'h058d: q1 = 16'h4a5f; // 0x0b1a
	13'h058e: q1 = 16'h226d; // 0x0b1c
	13'h058f: q1 = 16'h0024; // 0x0b1e
	13'h0590: q1 = 16'hd051; // 0x0b20
	13'h0591: q1 = 16'h3e00; // 0x0b22
	13'h0592: q1 = 16'hbe7c; // 0x0b24
	13'h0593: q1 = 16'h0280; // 0x0b26
	13'h0594: q1 = 16'h6c06; // 0x0b28
	13'h0595: q1 = 16'h3e3c; // 0x0b2a
	13'h0596: q1 = 16'h0280; // 0x0b2c
	13'h0597: q1 = 16'h600a; // 0x0b2e
	13'h0598: q1 = 16'hbe7c; // 0x0b30
	13'h0599: q1 = 16'h7580; // 0x0b32
	13'h059a: q1 = 16'h6d04; // 0x0b34
	13'h059b: q1 = 16'h3e3c; // 0x0b36
	13'h059c: q1 = 16'h7580; // 0x0b38
	13'h059d: q1 = 16'h206d; // 0x0b3a
	13'h059e: q1 = 16'h0024; // 0x0b3c
	13'h059f: q1 = 16'h3010; // 0x0b3e
	13'h05a0: q1 = 16'hb047; // 0x0b40
	13'h05a1: q1 = 16'h6606; // 0x0b42
	13'h05a2: q1 = 16'h3d7c; // 0x0b44
	13'h05a3: q1 = 16'h0001; // 0x0b46
	13'h05a4: q1 = 16'hfffe; // 0x0b48
	13'h05a5: q1 = 16'h206d; // 0x0b4a
	13'h05a6: q1 = 16'h0024; // 0x0b4c
	13'h05a7: q1 = 16'h3087; // 0x0b4e
	13'h05a8: q1 = 16'h206d; // 0x0b50
	13'h05a9: q1 = 16'h0020; // 0x0b52
	13'h05aa: q1 = 16'h3087; // 0x0b54
	13'h05ab: q1 = 16'h206d; // 0x0b56
	13'h05ac: q1 = 16'h002c; // 0x0b58
	13'h05ad: q1 = 16'h3087; // 0x0b5a
	13'h05ae: q1 = 16'h3ead; // 0x0b5c
	13'h05af: q1 = 16'h0010; // 0x0b5e
	13'h05b0: q1 = 16'h3f2d; // 0x0b60
	13'h05b1: q1 = 16'h000e; // 0x0b62
	13'h05b2: q1 = 16'h4eb9; // 0x0b64
	13'h05b3: q1 = 16'h0000; // 0x0b66
	13'h05b4: q1 = 16'ha730; // 0x0b68
	13'h05b5: q1 = 16'h4a5f; // 0x0b6a
	13'h05b6: q1 = 16'h3e00; // 0x0b6c
	13'h05b7: q1 = 16'hde6d; // 0x0b6e
	13'h05b8: q1 = 16'h0030; // 0x0b70
	13'h05b9: q1 = 16'hbe7c; // 0x0b72
	13'h05ba: q1 = 16'h1500; // 0x0b74
	13'h05bb: q1 = 16'h6c06; // 0x0b76
	13'h05bc: q1 = 16'h3e3c; // 0x0b78
	13'h05bd: q1 = 16'h1500; // 0x0b7a
	13'h05be: q1 = 16'h600a; // 0x0b7c
	13'h05bf: q1 = 16'hbe7c; // 0x0b7e
	13'h05c0: q1 = 16'h7400; // 0x0b80
	13'h05c1: q1 = 16'h6d04; // 0x0b82
	13'h05c2: q1 = 16'h3e3c; // 0x0b84
	13'h05c3: q1 = 16'h7400; // 0x0b86
	13'h05c4: q1 = 16'hbe6d; // 0x0b88
	13'h05c5: q1 = 16'h0030; // 0x0b8a
	13'h05c6: q1 = 16'h6606; // 0x0b8c
	13'h05c7: q1 = 16'h3d7c; // 0x0b8e
	13'h05c8: q1 = 16'h0001; // 0x0b90
	13'h05c9: q1 = 16'hfffc; // 0x0b92
	13'h05ca: q1 = 16'h4a6e; // 0x0b94
	13'h05cb: q1 = 16'hfffe; // 0x0b96
	13'h05cc: q1 = 16'h670a; // 0x0b98
	13'h05cd: q1 = 16'h4a6e; // 0x0b9a
	13'h05ce: q1 = 16'hfffc; // 0x0b9c
	13'h05cf: q1 = 16'h6704; // 0x0b9e
	13'h05d0: q1 = 16'h426d; // 0x0ba0
	13'h05d1: q1 = 16'h0010; // 0x0ba2
	13'h05d2: q1 = 16'h3c15; // 0x0ba4
	13'h05d3: q1 = 16'h3b47; // 0x0ba6
	13'h05d4: q1 = 16'h0030; // 0x0ba8
	13'h05d5: q1 = 16'h4a6d; // 0x0baa
	13'h05d6: q1 = 16'h0010; // 0x0bac
	13'h05d7: q1 = 16'h6f0e; // 0x0bae
	13'h05d8: q1 = 16'h4a46; // 0x0bb0
	13'h05d9: q1 = 16'h6706; // 0x0bb2
	13'h05da: q1 = 16'hbc7c; // 0x0bb4
	13'h05db: q1 = 16'h0004; // 0x0bb6
	13'h05dc: q1 = 16'h6604; // 0x0bb8
	13'h05dd: q1 = 16'hde7c; // 0x0bba
	13'h05de: q1 = 16'h0080; // 0x0bbc
	13'h05df: q1 = 16'h206d; // 0x0bbe
	13'h05e0: q1 = 16'h0024; // 0x0bc0
	13'h05e1: q1 = 16'h3147; // 0x0bc2
	13'h05e2: q1 = 16'h0002; // 0x0bc4
	13'h05e3: q1 = 16'h206d; // 0x0bc6
	13'h05e4: q1 = 16'h0020; // 0x0bc8
	13'h05e5: q1 = 16'h3207; // 0x0bca
	13'h05e6: q1 = 16'hd27c; // 0x0bcc
	13'h05e7: q1 = 16'h0200; // 0x0bce
	13'h05e8: q1 = 16'h3141; // 0x0bd0
	13'h05e9: q1 = 16'h0002; // 0x0bd2
	13'h05ea: q1 = 16'h206d; // 0x0bd4
	13'h05eb: q1 = 16'h002c; // 0x0bd6
	13'h05ec: q1 = 16'h226d; // 0x0bd8
	13'h05ed: q1 = 16'h0020; // 0x0bda
	13'h05ee: q1 = 16'h3169; // 0x0bdc
	13'h05ef: q1 = 16'h0002; // 0x0bde
	13'h05f0: q1 = 16'h0002; // 0x0be0
	13'h05f1: q1 = 16'h4a6d; // 0x0be2
	13'h05f2: q1 = 16'h0010; // 0x0be4
	13'h05f3: q1 = 16'h673c; // 0x0be6
	13'h05f4: q1 = 16'h4a6d; // 0x0be8
	13'h05f5: q1 = 16'h0002; // 0x0bea
	13'h05f6: q1 = 16'h6632; // 0x0bec
	13'h05f7: q1 = 16'h3b6d; // 0x0bee
	13'h05f8: q1 = 16'h0004; // 0x0bf0
	13'h05f9: q1 = 16'h0002; // 0x0bf2
	13'h05fa: q1 = 16'h5255; // 0x0bf4
	13'h05fb: q1 = 16'h0c55; // 0x0bf6
	13'h05fc: q1 = 16'h0008; // 0x0bf8
	13'h05fd: q1 = 16'h6602; // 0x0bfa
	13'h05fe: q1 = 16'h4255; // 0x0bfc
	13'h05ff: q1 = 16'h0c55; // 0x0bfe
	13'h0600: q1 = 16'h0002; // 0x0c00
	13'h0601: q1 = 16'h6706; // 0x0c02
	13'h0602: q1 = 16'h0c55; // 0x0c04
	13'h0603: q1 = 16'h0006; // 0x0c06
	13'h0604: q1 = 16'h6614; // 0x0c08
	13'h0605: q1 = 16'h4a79; // 0x0c0a
	13'h0606: q1 = 16'h0001; // 0x0c0c
	13'h0607: q1 = 16'h8676; // 0x0c0e
	13'h0608: q1 = 16'h660c; // 0x0c10
	13'h0609: q1 = 16'h2ebc; // 0x0c12
	13'h060a: q1 = 16'h0000; // 0x0c14
	13'h060b: q1 = 16'hfd1c; // 0x0c16
	13'h060c: q1 = 16'h4eb9; // 0x0c18
	13'h060d: q1 = 16'h0000; // 0x0c1a
	13'h060e: q1 = 16'h7dd8; // 0x0c1c
	13'h060f: q1 = 16'h6004; // 0x0c1e
	13'h0610: q1 = 16'h536d; // 0x0c20
	13'h0611: q1 = 16'h0002; // 0x0c22
	13'h0612: q1 = 16'h4a6d; // 0x0c24
	13'h0613: q1 = 16'h0010; // 0x0c26
	13'h0614: q1 = 16'h671a; // 0x0c28
	13'h0615: q1 = 16'h206d; // 0x0c2a
	13'h0616: q1 = 16'h0024; // 0x0c2c
	13'h0617: q1 = 16'h3215; // 0x0c2e
	13'h0618: q1 = 16'h48c1; // 0x0c30
	13'h0619: q1 = 16'hd2bc; // 0x0c32
	13'h061a: q1 = 16'h0000; // 0x0c34
	13'h061b: q1 = 16'hcb5a; // 0x0c36
	13'h061c: q1 = 16'h2241; // 0x0c38
	13'h061d: q1 = 16'h1211; // 0x0c3a
	13'h061e: q1 = 16'h4881; // 0x0c3c
	13'h061f: q1 = 16'h3141; // 0x0c3e
	13'h0620: q1 = 16'h0004; // 0x0c40
	13'h0621: q1 = 16'h600a; // 0x0c42
	13'h0622: q1 = 16'h206d; // 0x0c44
	13'h0623: q1 = 16'h0024; // 0x0c46
	13'h0624: q1 = 16'h317c; // 0x0c48
	13'h0625: q1 = 16'h00bf; // 0x0c4a
	13'h0626: q1 = 16'h0004; // 0x0c4c
	13'h0627: q1 = 16'h302d; // 0x0c4e
	13'h0628: q1 = 16'h000e; // 0x0c50
	13'h0629: q1 = 16'h48c0; // 0x0c52
	13'h062a: q1 = 16'hd0bc; // 0x0c54
	13'h062b: q1 = 16'h0000; // 0x0c56
	13'h062c: q1 = 16'hca18; // 0x0c58
	13'h062d: q1 = 16'h2040; // 0x0c5a
	13'h062e: q1 = 16'h1e10; // 0x0c5c
	13'h062f: q1 = 16'h4887; // 0x0c5e
	13'h0630: q1 = 16'h4aad; // 0x0c60
	13'h0631: q1 = 16'h0006; // 0x0c62
	13'h0632: q1 = 16'h661a; // 0x0c64
	13'h0633: q1 = 16'h206d; // 0x0c66
	13'h0634: q1 = 16'h002c; // 0x0c68
	13'h0635: q1 = 16'h3207; // 0x0c6a
	13'h0636: q1 = 16'h48c1; // 0x0c6c
	13'h0637: q1 = 16'hd2bc; // 0x0c6e
	13'h0638: q1 = 16'h0000; // 0x0c70
	13'h0639: q1 = 16'hcb62; // 0x0c72
	13'h063a: q1 = 16'h2241; // 0x0c74
	13'h063b: q1 = 16'h1211; // 0x0c76
	13'h063c: q1 = 16'h4881; // 0x0c78
	13'h063d: q1 = 16'h3141; // 0x0c7a
	13'h063e: q1 = 16'h0004; // 0x0c7c
	13'h063f: q1 = 16'h600e; // 0x0c7e
	13'h0640: q1 = 16'h206d; // 0x0c80
	13'h0641: q1 = 16'h002c; // 0x0c82
	13'h0642: q1 = 16'h3207; // 0x0c84
	13'h0643: q1 = 16'hd27c; // 0x0c86
	13'h0644: q1 = 16'h00df; // 0x0c88
	13'h0645: q1 = 16'h3141; // 0x0c8a
	13'h0646: q1 = 16'h0004; // 0x0c8c
	13'h0647: q1 = 16'h206d; // 0x0c8e
	13'h0648: q1 = 16'h0020; // 0x0c90
	13'h0649: q1 = 16'h3207; // 0x0c92
	13'h064a: q1 = 16'hd27c; // 0x0c94
	13'h064b: q1 = 16'h000c; // 0x0c96
	13'h064c: q1 = 16'h3141; // 0x0c98
	13'h064d: q1 = 16'h0004; // 0x0c9a
	13'h064e: q1 = 16'h0c6d; // 0x0c9c
	13'h064f: q1 = 16'h0004; // 0x0c9e
	13'h0650: q1 = 16'h001a; // 0x0ca0
	13'h0651: q1 = 16'h6700; // 0x0ca2
	13'h0652: q1 = 16'h007a; // 0x0ca4
	13'h0653: q1 = 16'h4a6e; // 0x0ca6
	13'h0654: q1 = 16'hfff8; // 0x0ca8
	13'h0655: q1 = 16'h6742; // 0x0caa
	13'h0656: q1 = 16'h4aad; // 0x0cac
	13'h0657: q1 = 16'h0006; // 0x0cae
	13'h0658: q1 = 16'h673c; // 0x0cb0
	13'h0659: q1 = 16'h4aad; // 0x0cb2
	13'h065a: q1 = 16'h001c; // 0x0cb4
	13'h065b: q1 = 16'h6636; // 0x0cb6
	13'h065c: q1 = 16'h2b7c; // 0x0cb8
	13'h065d: q1 = 16'h0000; // 0x0cba
	13'h065e: q1 = 16'h0005; // 0x0cbc
	13'h065f: q1 = 16'h001c; // 0x0cbe
	13'h0660: q1 = 16'h2eb9; // 0x0cc0
	13'h0661: q1 = 16'h0000; // 0x0cc2
	13'h0662: q1 = 16'hcb06; // 0x0cc4
	13'h0663: q1 = 16'h3f2d; // 0x0cc6
	13'h0664: q1 = 16'h000e; // 0x0cc8
	13'h0665: q1 = 16'h2f2d; // 0x0cca
	13'h0666: q1 = 16'h0006; // 0x0ccc
	13'h0667: q1 = 16'h4eb9; // 0x0cce
	13'h0668: q1 = 16'h0000; // 0x0cd0
	13'h0669: q1 = 16'h3b8e; // 0x0cd2
	13'h066a: q1 = 16'h5c4f; // 0x0cd4
	13'h066b: q1 = 16'h4a79; // 0x0cd6
	13'h066c: q1 = 16'h0001; // 0x0cd8
	13'h066d: q1 = 16'h8676; // 0x0cda
	13'h066e: q1 = 16'h660c; // 0x0cdc
	13'h066f: q1 = 16'h2ebc; // 0x0cde
	13'h0670: q1 = 16'h0000; // 0x0ce0
	13'h0671: q1 = 16'hfdf8; // 0x0ce2
	13'h0672: q1 = 16'h4eb9; // 0x0ce4
	13'h0673: q1 = 16'h0000; // 0x0ce6
	13'h0674: q1 = 16'h7dd8; // 0x0ce8
	13'h0675: q1 = 16'h42ad; // 0x0cea
	13'h0676: q1 = 16'h0006; // 0x0cec
	13'h0677: q1 = 16'h4aad; // 0x0cee
	13'h0678: q1 = 16'h0006; // 0x0cf0
	13'h0679: q1 = 16'h662a; // 0x0cf2
	13'h067a: q1 = 16'h202d; // 0x0cf4
	13'h067b: q1 = 16'h001c; // 0x0cf6
	13'h067c: q1 = 16'h4a40; // 0x0cf8
	13'h067d: q1 = 16'h6704; // 0x0cfa
	13'h067e: q1 = 16'h4257; // 0x0cfc
	13'h067f: q1 = 16'h6004; // 0x0cfe
	13'h0680: q1 = 16'h3ebc; // 0x0d00
	13'h0681: q1 = 16'h0001; // 0x0d02
	13'h0682: q1 = 16'h206d; // 0x0d04
	13'h0683: q1 = 16'h0024; // 0x0d06
	13'h0684: q1 = 16'h3f28; // 0x0d08
	13'h0685: q1 = 16'h0002; // 0x0d0a
	13'h0686: q1 = 16'h206d; // 0x0d0c
	13'h0687: q1 = 16'h0024; // 0x0d0e
	13'h0688: q1 = 16'h3f10; // 0x0d10
	13'h0689: q1 = 16'h4eb9; // 0x0d12
	13'h068a: q1 = 16'h0000; // 0x0d14
	13'h068b: q1 = 16'h37e6; // 0x0d16
	13'h068c: q1 = 16'h4a9f; // 0x0d18
	13'h068d: q1 = 16'h2b40; // 0x0d1a
	13'h068e: q1 = 16'h0006; // 0x0d1c
	13'h068f: q1 = 16'h4eb9; // 0x0d1e
	13'h0690: q1 = 16'h0000; // 0x0d20
	13'h0691: q1 = 16'h607a; // 0x0d22
	13'h0692: q1 = 16'h3ead; // 0x0d24
	13'h0693: q1 = 16'h000e; // 0x0d26
	13'h0694: q1 = 16'h202d; // 0x0d28
	13'h0695: q1 = 16'h0024; // 0x0d2a
	13'h0696: q1 = 16'h5c80; // 0x0d2c
	13'h0697: q1 = 16'h2f00; // 0x0d2e
	13'h0698: q1 = 16'h4eb9; // 0x0d30
	13'h0699: q1 = 16'h0000; // 0x0d32
	13'h069a: q1 = 16'h3ee6; // 0x0d34
	13'h069b: q1 = 16'h4a9f; // 0x0d36
	13'h069c: q1 = 16'h3ead; // 0x0d38
	13'h069d: q1 = 16'h000e; // 0x0d3a
	13'h069e: q1 = 16'h202d; // 0x0d3c
	13'h069f: q1 = 16'h0028; // 0x0d3e
	13'h06a0: q1 = 16'h5c80; // 0x0d40
	13'h06a1: q1 = 16'h2f00; // 0x0d42
	13'h06a2: q1 = 16'h4eb9; // 0x0d44
	13'h06a3: q1 = 16'h0000; // 0x0d46
	13'h06a4: q1 = 16'h3ee6; // 0x0d48
	13'h06a5: q1 = 16'h4a9f; // 0x0d4a
	13'h06a6: q1 = 16'h3ead; // 0x0d4c
	13'h06a7: q1 = 16'h000e; // 0x0d4e
	13'h06a8: q1 = 16'h202d; // 0x0d50
	13'h06a9: q1 = 16'h0020; // 0x0d52
	13'h06aa: q1 = 16'h5c80; // 0x0d54
	13'h06ab: q1 = 16'h2f00; // 0x0d56
	13'h06ac: q1 = 16'h4eb9; // 0x0d58
	13'h06ad: q1 = 16'h0000; // 0x0d5a
	13'h06ae: q1 = 16'h3ee6; // 0x0d5c
	13'h06af: q1 = 16'h4a9f; // 0x0d5e
	13'h06b0: q1 = 16'h3ead; // 0x0d60
	13'h06b1: q1 = 16'h000e; // 0x0d62
	13'h06b2: q1 = 16'h202d; // 0x0d64
	13'h06b3: q1 = 16'h002c; // 0x0d66
	13'h06b4: q1 = 16'h5c80; // 0x0d68
	13'h06b5: q1 = 16'h2f00; // 0x0d6a
	13'h06b6: q1 = 16'h4eb9; // 0x0d6c
	13'h06b7: q1 = 16'h0000; // 0x0d6e
	13'h06b8: q1 = 16'h3ee6; // 0x0d70
	13'h06b9: q1 = 16'h4a9f; // 0x0d72
	13'h06ba: q1 = 16'h4a9f; // 0x0d74
	13'h06bb: q1 = 16'h4cdf; // 0x0d76
	13'h06bc: q1 = 16'h38f8; // 0x0d78
	13'h06bd: q1 = 16'h4e5e; // 0x0d7a
	13'h06be: q1 = 16'h4e75; // 0x0d7c
	13'h06bf: q1 = 16'h4e56; // 0x0d7e
	13'h06c0: q1 = 16'hfffe; // 0x0d80
	13'h06c1: q1 = 16'h48e7; // 0x0d82
	13'h06c2: q1 = 16'h0104; // 0x0d84
	13'h06c3: q1 = 16'h2a7c; // 0x0d86
	13'h06c4: q1 = 16'h0001; // 0x0d88
	13'h06c5: q1 = 16'h7f2c; // 0x0d8a
	13'h06c6: q1 = 16'h206d; // 0x0d8c
	13'h06c7: q1 = 16'h0024; // 0x0d8e
	13'h06c8: q1 = 16'h3010; // 0x0d90
	13'h06c9: q1 = 16'h906e; // 0x0d92
	13'h06ca: q1 = 16'h0008; // 0x0d94
	13'h06cb: q1 = 16'h3d40; // 0x0d96
	13'h06cc: q1 = 16'hfffe; // 0x0d98
	13'h06cd: q1 = 16'h4a6e; // 0x0d9a
	13'h06ce: q1 = 16'hfffe; // 0x0d9c
	13'h06cf: q1 = 16'h6c0a; // 0x0d9e
	13'h06d0: q1 = 16'h302e; // 0x0da0
	13'h06d1: q1 = 16'hfffe; // 0x0da2
	13'h06d2: q1 = 16'h4440; // 0x0da4
	13'h06d3: q1 = 16'h3d40; // 0x0da6
	13'h06d4: q1 = 16'hfffe; // 0x0da8
	13'h06d5: q1 = 16'h0c6e; // 0x0daa
	13'h06d6: q1 = 16'h1800; // 0x0dac
	13'h06d7: q1 = 16'hfffe; // 0x0dae
	13'h06d8: q1 = 16'h6f04; // 0x0db0
	13'h06d9: q1 = 16'h4240; // 0x0db2
	13'h06da: q1 = 16'h602e; // 0x0db4
	13'h06db: q1 = 16'h206d; // 0x0db6
	13'h06dc: q1 = 16'h0024; // 0x0db8
	13'h06dd: q1 = 16'h3028; // 0x0dba
	13'h06de: q1 = 16'h0002; // 0x0dbc
	13'h06df: q1 = 16'h906e; // 0x0dbe
	13'h06e0: q1 = 16'h000a; // 0x0dc0
	13'h06e1: q1 = 16'h3d40; // 0x0dc2
	13'h06e2: q1 = 16'hfffe; // 0x0dc4
	13'h06e3: q1 = 16'h4a6e; // 0x0dc6
	13'h06e4: q1 = 16'hfffe; // 0x0dc8
	13'h06e5: q1 = 16'h6c0a; // 0x0dca
	13'h06e6: q1 = 16'h302e; // 0x0dcc
	13'h06e7: q1 = 16'hfffe; // 0x0dce
	13'h06e8: q1 = 16'h4440; // 0x0dd0
	13'h06e9: q1 = 16'h3d40; // 0x0dd2
	13'h06ea: q1 = 16'hfffe; // 0x0dd4
	13'h06eb: q1 = 16'h0c6e; // 0x0dd6
	13'h06ec: q1 = 16'h1800; // 0x0dd8
	13'h06ed: q1 = 16'hfffe; // 0x0dda
	13'h06ee: q1 = 16'h6f04; // 0x0ddc
	13'h06ef: q1 = 16'h4240; // 0x0dde
	13'h06f0: q1 = 16'h6002; // 0x0de0
	13'h06f1: q1 = 16'h7001; // 0x0de2
	13'h06f2: q1 = 16'h4a9f; // 0x0de4
	13'h06f3: q1 = 16'h4cdf; // 0x0de6
	13'h06f4: q1 = 16'h2000; // 0x0de8
	13'h06f5: q1 = 16'h4e5e; // 0x0dea
	13'h06f6: q1 = 16'h4e75; // 0x0dec
	13'h06f7: q1 = 16'h4e56; // 0x0dee
	13'h06f8: q1 = 16'h0000; // 0x0df0
	13'h06f9: q1 = 16'h48e7; // 0x0df2
	13'h06fa: q1 = 16'h0104; // 0x0df4
	13'h06fb: q1 = 16'h2a7c; // 0x0df6
	13'h06fc: q1 = 16'h0001; // 0x0df8
	13'h06fd: q1 = 16'h7f2c; // 0x0dfa
	13'h06fe: q1 = 16'h4a79; // 0x0dfc
	13'h06ff: q1 = 16'h0001; // 0x0dfe
	13'h0700: q1 = 16'h8676; // 0x0e00
	13'h0701: q1 = 16'h670a; // 0x0e02
	13'h0702: q1 = 16'h2b79; // 0x0e04
	13'h0703: q1 = 16'h0001; // 0x0e06
	13'h0704: q1 = 16'h7fb2; // 0x0e08
	13'h0705: q1 = 16'h0006; // 0x0e0a
	13'h0706: q1 = 16'h6008; // 0x0e0c
	13'h0707: q1 = 16'h23ed; // 0x0e0e
	13'h0708: q1 = 16'h0006; // 0x0e10
	13'h0709: q1 = 16'h0001; // 0x0e12
	13'h070a: q1 = 16'h7fb2; // 0x0e14
	13'h070b: q1 = 16'h206d; // 0x0e16
	13'h070c: q1 = 16'h0024; // 0x0e18
	13'h070d: q1 = 16'h30bc; // 0x0e1a
	13'h070e: q1 = 16'h7380; // 0x0e1c
	13'h070f: q1 = 16'h206d; // 0x0e1e
	13'h0710: q1 = 16'h0024; // 0x0e20
	13'h0711: q1 = 16'h323c; // 0x0e22
	13'h0712: q1 = 16'h1400; // 0x0e24
	13'h0713: q1 = 16'h9279; // 0x0e26
	13'h0714: q1 = 16'h0001; // 0x0e28
	13'h0715: q1 = 16'h8938; // 0x0e2a
	13'h0716: q1 = 16'hd27c; // 0x0e2c
	13'h0717: q1 = 16'h7400; // 0x0e2e
	13'h0718: q1 = 16'h3141; // 0x0e30
	13'h0719: q1 = 16'h0002; // 0x0e32
	13'h071a: q1 = 16'h4a79; // 0x0e34
	13'h071b: q1 = 16'h0001; // 0x0e36
	13'h071c: q1 = 16'h8676; // 0x0e38
	13'h071d: q1 = 16'h671a; // 0x0e3a
	13'h071e: q1 = 16'h2039; // 0x0e3c
	13'h071f: q1 = 16'h0001; // 0x0e3e
	13'h0720: q1 = 16'h86ae; // 0x0e40
	13'h0721: q1 = 16'h90bc; // 0x0e42
	13'h0722: q1 = 16'h0001; // 0x0e44
	13'h0723: q1 = 16'h81fe; // 0x0e46
	13'h0724: q1 = 16'hd0bc; // 0x0e48
	13'h0725: q1 = 16'h0000; // 0x0e4a
	13'h0726: q1 = 16'h0017; // 0x0e4c
	13'h0727: q1 = 16'h3e80; // 0x0e4e
	13'h0728: q1 = 16'h4eb9; // 0x0e50
	13'h0729: q1 = 16'h0000; // 0x0e52
	13'h072a: q1 = 16'h7d88; // 0x0e54
	13'h072b: q1 = 16'h23fc; // 0x0e56
	13'h072c: q1 = 16'h0001; // 0x0e58
	13'h072d: q1 = 16'h81fe; // 0x0e5a
	13'h072e: q1 = 16'h0001; // 0x0e5c
	13'h072f: q1 = 16'h86ae; // 0x0e5e
	13'h0730: q1 = 16'h23fc; // 0x0e60
	13'h0731: q1 = 16'h0001; // 0x0e62
	13'h0732: q1 = 16'h8882; // 0x0e64
	13'h0733: q1 = 16'h0001; // 0x0e66
	13'h0734: q1 = 16'h7ebc; // 0x0e68
	13'h0735: q1 = 16'h4279; // 0x0e6a
	13'h0736: q1 = 16'h0001; // 0x0e6c
	13'h0737: q1 = 16'h7ba2; // 0x0e6e
	13'h0738: q1 = 16'h4279; // 0x0e70
	13'h0739: q1 = 16'h0001; // 0x0e72
	13'h073a: q1 = 16'h7f22; // 0x0e74
	13'h073b: q1 = 16'h4279; // 0x0e76
	13'h073c: q1 = 16'h0001; // 0x0e78
	13'h073d: q1 = 16'h7efc; // 0x0e7a
	13'h073e: q1 = 16'h3b7c; // 0x0e7c
	13'h073f: q1 = 16'h0024; // 0x0e7e
	13'h0740: q1 = 16'h000e; // 0x0e80
	13'h0741: q1 = 16'h4eb9; // 0x0e82
	13'h0742: q1 = 16'h0000; // 0x0e84
	13'h0743: q1 = 16'h61f8; // 0x0e86
	13'h0744: q1 = 16'h4aad; // 0x0e88
	13'h0745: q1 = 16'h0006; // 0x0e8a
	13'h0746: q1 = 16'h671e; // 0x0e8c
	13'h0747: q1 = 16'h206d; // 0x0e8e
	13'h0748: q1 = 16'h002c; // 0x0e90
	13'h0749: q1 = 16'h322d; // 0x0e92
	13'h074a: q1 = 16'h000e; // 0x0e94
	13'h074b: q1 = 16'h48c1; // 0x0e96
	13'h074c: q1 = 16'hd2bc; // 0x0e98
	13'h074d: q1 = 16'h0000; // 0x0e9a
	13'h074e: q1 = 16'hca18; // 0x0e9c
	13'h074f: q1 = 16'h2241; // 0x0e9e
	13'h0750: q1 = 16'h1211; // 0x0ea0
	13'h0751: q1 = 16'h4881; // 0x0ea2
	13'h0752: q1 = 16'hd27c; // 0x0ea4
	13'h0753: q1 = 16'h00df; // 0x0ea6
	13'h0754: q1 = 16'h3141; // 0x0ea8
	13'h0755: q1 = 16'h0004; // 0x0eaa
	13'h0756: q1 = 16'h2ead; // 0x0eac
	13'h0757: q1 = 16'h0006; // 0x0eae
	13'h0758: q1 = 16'h4eb9; // 0x0eb0
	13'h0759: q1 = 16'h0000; // 0x0eb2
	13'h075a: q1 = 16'h3a7c; // 0x0eb4
	13'h075b: q1 = 16'h4eb9; // 0x0eb6
	13'h075c: q1 = 16'h0000; // 0x0eb8
	13'h075d: q1 = 16'h607a; // 0x0eba
	13'h075e: q1 = 16'h4a9f; // 0x0ebc
	13'h075f: q1 = 16'h4cdf; // 0x0ebe
	13'h0760: q1 = 16'h2000; // 0x0ec0
	13'h0761: q1 = 16'h4e5e; // 0x0ec2
	13'h0762: q1 = 16'h4e75; // 0x0ec4
	13'h0763: q1 = 16'h4e56; // 0x0ec6
	13'h0764: q1 = 16'h0000; // 0x0ec8
	13'h0765: q1 = 16'h48e7; // 0x0eca
	13'h0766: q1 = 16'h0104; // 0x0ecc
	13'h0767: q1 = 16'h2a7c; // 0x0ece
	13'h0768: q1 = 16'h0001; // 0x0ed0
	13'h0769: q1 = 16'h7f2c; // 0x0ed2
	13'h076a: q1 = 16'h302d; // 0x0ed4
	13'h076b: q1 = 16'h001a; // 0x0ed6
	13'h076c: q1 = 16'h4a9f; // 0x0ed8
	13'h076d: q1 = 16'h4cdf; // 0x0eda
	13'h076e: q1 = 16'h2000; // 0x0edc
	13'h076f: q1 = 16'h4e5e; // 0x0ede
	13'h0770: q1 = 16'h4e75; // 0x0ee0
	13'h0771: q1 = 16'h4e56; // 0x0ee2
	13'h0772: q1 = 16'h0000; // 0x0ee4
	13'h0773: q1 = 16'h48e7; // 0x0ee6
	13'h0774: q1 = 16'h0104; // 0x0ee8
	13'h0775: q1 = 16'h2a7c; // 0x0eea
	13'h0776: q1 = 16'h0001; // 0x0eec
	13'h0777: q1 = 16'h7f2c; // 0x0eee
	13'h0778: q1 = 16'h206d; // 0x0ef0
	13'h0779: q1 = 16'h0024; // 0x0ef2
	13'h077a: q1 = 16'h3010; // 0x0ef4
	13'h077b: q1 = 16'h4a9f; // 0x0ef6
	13'h077c: q1 = 16'h4cdf; // 0x0ef8
	13'h077d: q1 = 16'h2000; // 0x0efa
	13'h077e: q1 = 16'h4e5e; // 0x0efc
	13'h077f: q1 = 16'h4e75; // 0x0efe
	13'h0780: q1 = 16'h4e56; // 0x0f00
	13'h0781: q1 = 16'hfffe; // 0x0f02
	13'h0782: q1 = 16'h48e7; // 0x0f04
	13'h0783: q1 = 16'h0104; // 0x0f06
	13'h0784: q1 = 16'h2a7c; // 0x0f08
	13'h0785: q1 = 16'h0001; // 0x0f0a
	13'h0786: q1 = 16'h7f2c; // 0x0f0c
	13'h0787: q1 = 16'h3ead; // 0x0f0e
	13'h0788: q1 = 16'h0010; // 0x0f10
	13'h0789: q1 = 16'h3f2d; // 0x0f12
	13'h078a: q1 = 16'h000e; // 0x0f14
	13'h078b: q1 = 16'h4eb9; // 0x0f16
	13'h078c: q1 = 16'h0000; // 0x0f18
	13'h078d: q1 = 16'h1280; // 0x0f1a
	13'h078e: q1 = 16'h4a5f; // 0x0f1c
	13'h078f: q1 = 16'h3d40; // 0x0f1e
	13'h0790: q1 = 16'hfffe; // 0x0f20
	13'h0791: q1 = 16'h302e; // 0x0f22
	13'h0792: q1 = 16'hfffe; // 0x0f24
	13'h0793: q1 = 16'h4a9f; // 0x0f26
	13'h0794: q1 = 16'h4cdf; // 0x0f28
	13'h0795: q1 = 16'h2000; // 0x0f2a
	13'h0796: q1 = 16'h4e5e; // 0x0f2c
	13'h0797: q1 = 16'h4e75; // 0x0f2e
	13'h0798: q1 = 16'h4e56; // 0x0f30
	13'h0799: q1 = 16'h0000; // 0x0f32
	13'h079a: q1 = 16'h48e7; // 0x0f34
	13'h079b: q1 = 16'h0104; // 0x0f36
	13'h079c: q1 = 16'h2a7c; // 0x0f38
	13'h079d: q1 = 16'h0001; // 0x0f3a
	13'h079e: q1 = 16'h7f2c; // 0x0f3c
	13'h079f: q1 = 16'h206d; // 0x0f3e
	13'h07a0: q1 = 16'h0024; // 0x0f40
	13'h07a1: q1 = 16'h3028; // 0x0f42
	13'h07a2: q1 = 16'h0002; // 0x0f44
	13'h07a3: q1 = 16'h4a9f; // 0x0f46
	13'h07a4: q1 = 16'h4cdf; // 0x0f48
	13'h07a5: q1 = 16'h2000; // 0x0f4a
	13'h07a6: q1 = 16'h4e5e; // 0x0f4c
	13'h07a7: q1 = 16'h4e75; // 0x0f4e
	13'h07a8: q1 = 16'h4e56; // 0x0f50
	13'h07a9: q1 = 16'hfffe; // 0x0f52
	13'h07aa: q1 = 16'h48e7; // 0x0f54
	13'h07ab: q1 = 16'h0104; // 0x0f56
	13'h07ac: q1 = 16'h2a7c; // 0x0f58
	13'h07ad: q1 = 16'h0001; // 0x0f5a
	13'h07ae: q1 = 16'h7f2c; // 0x0f5c
	13'h07af: q1 = 16'h3ead; // 0x0f5e
	13'h07b0: q1 = 16'h0010; // 0x0f60
	13'h07b1: q1 = 16'h3f2d; // 0x0f62
	13'h07b2: q1 = 16'h000e; // 0x0f64
	13'h07b3: q1 = 16'h4eb9; // 0x0f66
	13'h07b4: q1 = 16'h0000; // 0x0f68
	13'h07b5: q1 = 16'ha730; // 0x0f6a
	13'h07b6: q1 = 16'h4a5f; // 0x0f6c
	13'h07b7: q1 = 16'h3d40; // 0x0f6e
	13'h07b8: q1 = 16'hfffe; // 0x0f70
	13'h07b9: q1 = 16'h302e; // 0x0f72
	13'h07ba: q1 = 16'hfffe; // 0x0f74
	13'h07bb: q1 = 16'h4a9f; // 0x0f76
	13'h07bc: q1 = 16'h4cdf; // 0x0f78
	13'h07bd: q1 = 16'h2000; // 0x0f7a
	13'h07be: q1 = 16'h4e5e; // 0x0f7c
	13'h07bf: q1 = 16'h4e75; // 0x0f7e
	13'h07c0: q1 = 16'h4e56; // 0x0f80
	13'h07c1: q1 = 16'hfff2; // 0x0f82
	13'h07c2: q1 = 16'h48e7; // 0x0f84
	13'h07c3: q1 = 16'h070c; // 0x0f86
	13'h07c4: q1 = 16'h2a7c; // 0x0f88
	13'h07c5: q1 = 16'h0001; // 0x0f8a
	13'h07c6: q1 = 16'h7f2c; // 0x0f8c
	13'h07c7: q1 = 16'h200e; // 0x0f8e
	13'h07c8: q1 = 16'hd0bc; // 0x0f90
	13'h07c9: q1 = 16'hffff; // 0x0f92
	13'h07ca: q1 = 16'hfff8; // 0x0f94
	13'h07cb: q1 = 16'h2e80; // 0x0f96
	13'h07cc: q1 = 16'h200e; // 0x0f98
	13'h07cd: q1 = 16'hd0bc; // 0x0f9a
	13'h07ce: q1 = 16'hffff; // 0x0f9c
	13'h07cf: q1 = 16'hfffa; // 0x0f9e
	13'h07d0: q1 = 16'h2f00; // 0x0fa0
	13'h07d1: q1 = 16'h200e; // 0x0fa2
	13'h07d2: q1 = 16'hd0bc; // 0x0fa4
	13'h07d3: q1 = 16'hffff; // 0x0fa6
	13'h07d4: q1 = 16'hfffc; // 0x0fa8
	13'h07d5: q1 = 16'h2f00; // 0x0faa
	13'h07d6: q1 = 16'h200e; // 0x0fac
	13'h07d7: q1 = 16'hd0bc; // 0x0fae
	13'h07d8: q1 = 16'hffff; // 0x0fb0
	13'h07d9: q1 = 16'hfffe; // 0x0fb2
	13'h07da: q1 = 16'h2f00; // 0x0fb4
	13'h07db: q1 = 16'h2f39; // 0x0fb6
	13'h07dc: q1 = 16'h0000; // 0x0fb8
	13'h07dd: q1 = 16'hcb14; // 0x0fba
	13'h07de: q1 = 16'h206d; // 0x0fbc
	13'h07df: q1 = 16'h0024; // 0x0fbe
	13'h07e0: q1 = 16'h3f28; // 0x0fc0
	13'h07e1: q1 = 16'h0002; // 0x0fc2
	13'h07e2: q1 = 16'h0657; // 0x0fc4
	13'h07e3: q1 = 16'h0200; // 0x0fc6
	13'h07e4: q1 = 16'h206d; // 0x0fc8
	13'h07e5: q1 = 16'h0024; // 0x0fca
	13'h07e6: q1 = 16'h3f10; // 0x0fcc
	13'h07e7: q1 = 16'h4eb9; // 0x0fce
	13'h07e8: q1 = 16'h0000; // 0x0fd0
	13'h07e9: q1 = 16'h36d8; // 0x0fd2
	13'h07ea: q1 = 16'hdefc; // 0x0fd4
	13'h07eb: q1 = 16'h0014; // 0x0fd6
	13'h07ec: q1 = 16'h2840; // 0x0fd8
	13'h07ed: q1 = 16'h0c79; // 0x0fda
	13'h07ee: q1 = 16'h0001; // 0x0fdc
	13'h07ef: q1 = 16'h0001; // 0x0fde
	13'h07f0: q1 = 16'h757c; // 0x0fe0
	13'h07f1: q1 = 16'h663c; // 0x0fe2
	13'h07f2: q1 = 16'h4a79; // 0x0fe4
	13'h07f3: q1 = 16'h0001; // 0x0fe6
	13'h07f4: q1 = 16'h7faa; // 0x0fe8
	13'h07f5: q1 = 16'h6634; // 0x0fea
	13'h07f6: q1 = 16'h2d79; // 0x0fec
	13'h07f7: q1 = 16'h0000; // 0x0fee
	13'h07f8: q1 = 16'hcb18; // 0x0ff0
	13'h07f9: q1 = 16'hfff4; // 0x0ff2
	13'h07fa: q1 = 16'h2039; // 0x0ff4
	13'h07fb: q1 = 16'h0000; // 0x0ff6
	13'h07fc: q1 = 16'hcb1c; // 0x0ff8
	13'h07fd: q1 = 16'he280; // 0x0ffa
	13'h07fe: q1 = 16'he380; // 0x0ffc
	13'h07ff: q1 = 16'hd1ae; // 0x0ffe
	13'h0800: q1 = 16'hfff4; // 0x1000
	13'h0801: q1 = 16'h206e; // 0x1002
	13'h0802: q1 = 16'hfff4; // 0x1004
	13'h0803: q1 = 16'h3d50; // 0x1006
	13'h0804: q1 = 16'hfff2; // 0x1008
	13'h0805: q1 = 16'h046e; // 0x100a
	13'h0806: q1 = 16'h2040; // 0x100c
	13'h0807: q1 = 16'hfff2; // 0x100e
	13'h0808: q1 = 16'h0c6e; // 0x1010
	13'h0809: q1 = 16'h0901; // 0x1012
	13'h080a: q1 = 16'hfff2; // 0x1014
	13'h080b: q1 = 16'h6708; // 0x1016
	13'h080c: q1 = 16'h33fc; // 0x1018
	13'h080d: q1 = 16'h0002; // 0x101a
	13'h080e: q1 = 16'h0001; // 0x101c
	13'h080f: q1 = 16'h757c; // 0x101e
	13'h0810: q1 = 16'h200c; // 0x1020
	13'h0811: q1 = 16'h675a; // 0x1022
	13'h0812: q1 = 16'h2e8c; // 0x1024
	13'h0813: q1 = 16'h4eb9; // 0x1026
	13'h0814: q1 = 16'h0000; // 0x1028
	13'h0815: q1 = 16'h3b7c; // 0x102a
	13'h0816: q1 = 16'h2b4c; // 0x102c
	13'h0817: q1 = 16'h000a; // 0x102e
	13'h0818: q1 = 16'h206d; // 0x1030
	13'h0819: q1 = 16'h0024; // 0x1032
	13'h081a: q1 = 16'h322e; // 0x1034
	13'h081b: q1 = 16'hfffe; // 0x1036
	13'h081c: q1 = 16'h5341; // 0x1038
	13'h081d: q1 = 16'he341; // 0x103a
	13'h081e: q1 = 16'h48c1; // 0x103c
	13'h081f: q1 = 16'hd2bc; // 0x103e
	13'h0820: q1 = 16'h0000; // 0x1040
	13'h0821: q1 = 16'hcb0a; // 0x1042
	13'h0822: q1 = 16'h2241; // 0x1044
	13'h0823: q1 = 16'h3151; // 0x1046
	13'h0824: q1 = 16'h0006; // 0x1048
	13'h0825: q1 = 16'h3b7c; // 0x104a
	13'h0826: q1 = 16'h0003; // 0x104c
	13'h0827: q1 = 16'h001a; // 0x104e
	13'h0828: q1 = 16'h206d; // 0x1050
	13'h0829: q1 = 16'h0024; // 0x1052
	13'h082a: q1 = 16'h317c; // 0x1054
	13'h082b: q1 = 16'h00bf; // 0x1056
	13'h082c: q1 = 16'h0004; // 0x1058
	13'h082d: q1 = 16'h206d; // 0x105a
	13'h082e: q1 = 16'h0028; // 0x105c
	13'h082f: q1 = 16'h317c; // 0x105e
	13'h0830: q1 = 16'h00be; // 0x1060
	13'h0831: q1 = 16'h0004; // 0x1062
	13'h0832: q1 = 16'h206d; // 0x1064
	13'h0833: q1 = 16'h0020; // 0x1066
	13'h0834: q1 = 16'h317c; // 0x1068
	13'h0835: q1 = 16'h008c; // 0x106a
	13'h0836: q1 = 16'h0004; // 0x106c
	13'h0837: q1 = 16'h206d; // 0x106e
	13'h0838: q1 = 16'h002c; // 0x1070
	13'h0839: q1 = 16'h317c; // 0x1072
	13'h083a: q1 = 16'h00cc; // 0x1074
	13'h083b: q1 = 16'h0004; // 0x1076
	13'h083c: q1 = 16'h7e01; // 0x1078
	13'h083d: q1 = 16'h6000; // 0x107a
	13'h083e: q1 = 16'h0134; // 0x107c
	13'h083f: q1 = 16'h4aad; // 0x107e
	13'h0840: q1 = 16'h001c; // 0x1080
	13'h0841: q1 = 16'h6622; // 0x1082
	13'h0842: q1 = 16'h3ead; // 0x1084
	13'h0843: q1 = 16'h0030; // 0x1086
	13'h0844: q1 = 16'h206d; // 0x1088
	13'h0845: q1 = 16'h0024; // 0x108a
	13'h0846: q1 = 16'h3f10; // 0x108c
	13'h0847: q1 = 16'h4eb9; // 0x108e
	13'h0848: q1 = 16'h0000; // 0x1090
	13'h0849: q1 = 16'h1e04; // 0x1092
	13'h084a: q1 = 16'h4a5f; // 0x1094
	13'h084b: q1 = 16'h4a40; // 0x1096
	13'h084c: q1 = 16'h670c; // 0x1098
	13'h084d: q1 = 16'h3b7c; // 0x109a
	13'h084e: q1 = 16'h0002; // 0x109c
	13'h084f: q1 = 16'h001a; // 0x109e
	13'h0850: q1 = 16'h7e01; // 0x10a0
	13'h0851: q1 = 16'h6000; // 0x10a2
	13'h0852: q1 = 16'h010c; // 0x10a4
	13'h0853: q1 = 16'h4eb9; // 0x10a6
	13'h0854: q1 = 16'h0000; // 0x10a8
	13'h0855: q1 = 16'h907c; // 0x10aa
	13'h0856: q1 = 16'h4a40; // 0x10ac
	13'h0857: q1 = 16'h6712; // 0x10ae
	13'h0858: q1 = 16'h3b7c; // 0x10b0
	13'h0859: q1 = 16'h0004; // 0x10b2
	13'h085a: q1 = 16'h001a; // 0x10b4
	13'h085b: q1 = 16'h3b7c; // 0x10b6
	13'h085c: q1 = 16'h00bc; // 0x10b8
	13'h085d: q1 = 16'h0010; // 0x10ba
	13'h085e: q1 = 16'h4247; // 0x10bc
	13'h085f: q1 = 16'h6000; // 0x10be
	13'h0860: q1 = 16'h00f0; // 0x10c0
	13'h0861: q1 = 16'h206d; // 0x10c2
	13'h0862: q1 = 16'h0024; // 0x10c4
	13'h0863: q1 = 16'h3d50; // 0x10c6
	13'h0864: q1 = 16'hfffa; // 0x10c8
	13'h0865: q1 = 16'h3d6d; // 0x10ca
	13'h0866: q1 = 16'h0030; // 0x10cc
	13'h0867: q1 = 16'hfff8; // 0x10ce
	13'h0868: q1 = 16'h4257; // 0x10d0
	13'h0869: q1 = 16'h200e; // 0x10d2
	13'h086a: q1 = 16'hd0bc; // 0x10d4
	13'h086b: q1 = 16'hffff; // 0x10d6
	13'h086c: q1 = 16'hfff8; // 0x10d8
	13'h086d: q1 = 16'h2f00; // 0x10da
	13'h086e: q1 = 16'h200e; // 0x10dc
	13'h086f: q1 = 16'hd0bc; // 0x10de
	13'h0870: q1 = 16'hffff; // 0x10e0
	13'h0871: q1 = 16'hfffa; // 0x10e2
	13'h0872: q1 = 16'h2f00; // 0x10e4
	13'h0873: q1 = 16'h4eb9; // 0x10e6
	13'h0874: q1 = 16'h0000; // 0x10e8
	13'h0875: q1 = 16'h5d44; // 0x10ea
	13'h0876: q1 = 16'hbf8f; // 0x10ec
	13'h0877: q1 = 16'h4a40; // 0x10ee
	13'h0878: q1 = 16'h6700; // 0x10f0
	13'h0879: q1 = 16'h00b8; // 0x10f2
	13'h087a: q1 = 16'h206d; // 0x10f4
	13'h087b: q1 = 16'h0024; // 0x10f6
	13'h087c: q1 = 16'h30ae; // 0x10f8
	13'h087d: q1 = 16'hfffa; // 0x10fa
	13'h087e: q1 = 16'h206d; // 0x10fc
	13'h087f: q1 = 16'h0024; // 0x10fe
	13'h0880: q1 = 16'h316e; // 0x1100
	13'h0881: q1 = 16'hfff8; // 0x1102
	13'h0882: q1 = 16'h0002; // 0x1104
	13'h0883: q1 = 16'h206d; // 0x1106
	13'h0884: q1 = 16'h0024; // 0x1108
	13'h0885: q1 = 16'h1239; // 0x110a
	13'h0886: q1 = 16'h0000; // 0x110c
	13'h0887: q1 = 16'hcb22; // 0x110e
	13'h0888: q1 = 16'h4881; // 0x1110
	13'h0889: q1 = 16'h3141; // 0x1112
	13'h088a: q1 = 16'h0004; // 0x1114
	13'h088b: q1 = 16'h206d; // 0x1116
	13'h088c: q1 = 16'h0028; // 0x1118
	13'h088d: q1 = 16'h30ae; // 0x111a
	13'h088e: q1 = 16'hfffa; // 0x111c
	13'h088f: q1 = 16'h206d; // 0x111e
	13'h0890: q1 = 16'h0028; // 0x1120
	13'h0891: q1 = 16'h316e; // 0x1122
	13'h0892: q1 = 16'hfff8; // 0x1124
	13'h0893: q1 = 16'h0002; // 0x1126
	13'h0894: q1 = 16'h206d; // 0x1128
	13'h0895: q1 = 16'h0028; // 0x112a
	13'h0896: q1 = 16'h1239; // 0x112c
	13'h0897: q1 = 16'h0000; // 0x112e
	13'h0898: q1 = 16'hcb46; // 0x1130
	13'h0899: q1 = 16'h4881; // 0x1132
	13'h089a: q1 = 16'h3141; // 0x1134
	13'h089b: q1 = 16'h0004; // 0x1136
	13'h089c: q1 = 16'h206d; // 0x1138
	13'h089d: q1 = 16'h0020; // 0x113a
	13'h089e: q1 = 16'h226d; // 0x113c
	13'h089f: q1 = 16'h0024; // 0x113e
	13'h08a0: q1 = 16'h3091; // 0x1140
	13'h08a1: q1 = 16'h206d; // 0x1142
	13'h08a2: q1 = 16'h0020; // 0x1144
	13'h08a3: q1 = 16'h226d; // 0x1146
	13'h08a4: q1 = 16'h0024; // 0x1148
	13'h08a5: q1 = 16'h3229; // 0x114a
	13'h08a6: q1 = 16'h0002; // 0x114c
	13'h08a7: q1 = 16'hd27c; // 0x114e
	13'h08a8: q1 = 16'h0200; // 0x1150
	13'h08a9: q1 = 16'h3141; // 0x1152
	13'h08aa: q1 = 16'h0002; // 0x1154
	13'h08ab: q1 = 16'h206d; // 0x1156
	13'h08ac: q1 = 16'h0020; // 0x1158
	13'h08ad: q1 = 16'h1239; // 0x115a
	13'h08ae: q1 = 16'h0000; // 0x115c
	13'h08af: q1 = 16'hcb2e; // 0x115e
	13'h08b0: q1 = 16'h4881; // 0x1160
	13'h08b1: q1 = 16'h3141; // 0x1162
	13'h08b2: q1 = 16'h0004; // 0x1164
	13'h08b3: q1 = 16'h206d; // 0x1166
	13'h08b4: q1 = 16'h002c; // 0x1168
	13'h08b5: q1 = 16'h226d; // 0x116a
	13'h08b6: q1 = 16'h0020; // 0x116c
	13'h08b7: q1 = 16'h3091; // 0x116e
	13'h08b8: q1 = 16'h206d; // 0x1170
	13'h08b9: q1 = 16'h002c; // 0x1172
	13'h08ba: q1 = 16'h226d; // 0x1174
	13'h08bb: q1 = 16'h0020; // 0x1176
	13'h08bc: q1 = 16'h3169; // 0x1178
	13'h08bd: q1 = 16'h0002; // 0x117a
	13'h08be: q1 = 16'h0002; // 0x117c
	13'h08bf: q1 = 16'h206d; // 0x117e
	13'h08c0: q1 = 16'h002c; // 0x1180
	13'h08c1: q1 = 16'h1239; // 0x1182
	13'h08c2: q1 = 16'h0000; // 0x1184
	13'h08c3: q1 = 16'hcb3a; // 0x1186
	13'h08c4: q1 = 16'h4881; // 0x1188
	13'h08c5: q1 = 16'h3141; // 0x118a
	13'h08c6: q1 = 16'h0004; // 0x118c
	13'h08c7: q1 = 16'h3b7c; // 0x118e
	13'h08c8: q1 = 16'h0001; // 0x1190
	13'h08c9: q1 = 16'h001a; // 0x1192
	13'h08ca: q1 = 16'h3b7c; // 0x1194
	13'h08cb: q1 = 16'h0002; // 0x1196
	13'h08cc: q1 = 16'h0012; // 0x1198
	13'h08cd: q1 = 16'h2ebc; // 0x119a
	13'h08ce: q1 = 16'h0000; // 0x119c
	13'h08cf: q1 = 16'hc972; // 0x119e
	13'h08d0: q1 = 16'h4eb9; // 0x11a0
	13'h08d1: q1 = 16'h0000; // 0x11a2
	13'h08d2: q1 = 16'h7dd8; // 0x11a4
	13'h08d3: q1 = 16'h7e01; // 0x11a6
	13'h08d4: q1 = 16'h6006; // 0x11a8
	13'h08d5: q1 = 16'h4240; // 0x11aa
	13'h08d6: q1 = 16'h6000; // 0x11ac
	13'h08d7: q1 = 16'h0092; // 0x11ae
	13'h08d8: q1 = 16'h4aad; // 0x11b0
	13'h08d9: q1 = 16'h0006; // 0x11b2
	13'h08da: q1 = 16'h670e; // 0x11b4
	13'h08db: q1 = 16'h2ead; // 0x11b6
	13'h08dc: q1 = 16'h0006; // 0x11b8
	13'h08dd: q1 = 16'h4eb9; // 0x11ba
	13'h08de: q1 = 16'h0000; // 0x11bc
	13'h08df: q1 = 16'h3356; // 0x11be
	13'h08e0: q1 = 16'h42ad; // 0x11c0
	13'h08e1: q1 = 16'h0006; // 0x11c2
	13'h08e2: q1 = 16'h4a47; // 0x11c4
	13'h08e3: q1 = 16'h6704; // 0x11c6
	13'h08e4: q1 = 16'h426d; // 0x11c8
	13'h08e5: q1 = 16'h0010; // 0x11ca
	13'h08e6: q1 = 16'h42ad; // 0x11cc
	13'h08e7: q1 = 16'h001c; // 0x11ce
	13'h08e8: q1 = 16'h4eb9; // 0x11d0
	13'h08e9: q1 = 16'h0000; // 0x11d2
	13'h08ea: q1 = 16'h607a; // 0x11d4
	13'h08eb: q1 = 16'h0c6d; // 0x11d6
	13'h08ec: q1 = 16'h0003; // 0x11d8
	13'h08ed: q1 = 16'h001a; // 0x11da
	13'h08ee: q1 = 16'h660e; // 0x11dc
	13'h08ef: q1 = 16'h206d; // 0x11de
	13'h08f0: q1 = 16'h0028; // 0x11e0
	13'h08f1: q1 = 16'h226d; // 0x11e2
	13'h08f2: q1 = 16'h0024; // 0x11e4
	13'h08f3: q1 = 16'h3169; // 0x11e6
	13'h08f4: q1 = 16'h0006; // 0x11e8
	13'h08f5: q1 = 16'h0006; // 0x11ea
	13'h08f6: q1 = 16'h4eb9; // 0x11ec
	13'h08f7: q1 = 16'h0000; // 0x11ee
	13'h08f8: q1 = 16'h90ec; // 0x11f0
	13'h08f9: q1 = 16'h3ebc; // 0x11f2
	13'h08fa: q1 = 16'h0001; // 0x11f4
	13'h08fb: q1 = 16'h4267; // 0x11f6
	13'h08fc: q1 = 16'h4eb9; // 0x11f8
	13'h08fd: q1 = 16'h0000; // 0x11fa
	13'h08fe: q1 = 16'h8e6c; // 0x11fc
	13'h08ff: q1 = 16'h4a5f; // 0x11fe
	13'h0900: q1 = 16'h3c00; // 0x1200
	13'h0901: q1 = 16'h2079; // 0x1202
	13'h0902: q1 = 16'h0001; // 0x1204
	13'h0903: q1 = 16'h7fb8; // 0x1206
	13'h0904: q1 = 16'h0c68; // 0x1208
	13'h0905: q1 = 16'h0001; // 0x120a
	13'h0906: q1 = 16'h0002; // 0x120c
	13'h0907: q1 = 16'h6602; // 0x120e
	13'h0908: q1 = 16'h7c01; // 0x1210
	13'h0909: q1 = 16'h0c6d; // 0x1212
	13'h090a: q1 = 16'h0001; // 0x1214
	13'h090b: q1 = 16'h001a; // 0x1216
	13'h090c: q1 = 16'h6724; // 0x1218
	13'h090d: q1 = 16'h3b7c; // 0x121a
	13'h090e: q1 = 16'h0001; // 0x121c
	13'h090f: q1 = 16'h0012; // 0x121e
	13'h0910: q1 = 16'h4a46; // 0x1220
	13'h0911: q1 = 16'h670e; // 0x1222
	13'h0912: q1 = 16'h2ebc; // 0x1224
	13'h0913: q1 = 16'h0000; // 0x1226
	13'h0914: q1 = 16'hc674; // 0x1228
	13'h0915: q1 = 16'h4eb9; // 0x122a
	13'h0916: q1 = 16'h0000; // 0x122c
	13'h0917: q1 = 16'h7ff8; // 0x122e
	13'h0918: q1 = 16'h600c; // 0x1230
	13'h0919: q1 = 16'h2ebc; // 0x1232
	13'h091a: q1 = 16'h0000; // 0x1234
	13'h091b: q1 = 16'hc6f2; // 0x1236
	13'h091c: q1 = 16'h4eb9; // 0x1238
	13'h091d: q1 = 16'h0000; // 0x123a
	13'h091e: q1 = 16'h7ff8; // 0x123c
	13'h091f: q1 = 16'h3007; // 0x123e
	13'h0920: q1 = 16'h4a9f; // 0x1240
	13'h0921: q1 = 16'h4cdf; // 0x1242
	13'h0922: q1 = 16'h30c0; // 0x1244
	13'h0923: q1 = 16'h4e5e; // 0x1246
	13'h0924: q1 = 16'h4e75; // 0x1248
	13'h0925: q1 = 16'h4e56; // 0x124a
	13'h0926: q1 = 16'h0000; // 0x124c
	13'h0927: q1 = 16'h48e7; // 0x124e
	13'h0928: q1 = 16'h0f04; // 0x1250
	13'h0929: q1 = 16'h2a7c; // 0x1252
	13'h092a: q1 = 16'h0001; // 0x1254
	13'h092b: q1 = 16'h7f2c; // 0x1256
	13'h092c: q1 = 16'h0c6d; // 0x1258
	13'h092d: q1 = 16'h0001; // 0x125a
	13'h092e: q1 = 16'h001a; // 0x125c
	13'h092f: q1 = 16'h6600; // 0x125e
	13'h0930: q1 = 16'h00e6; // 0x1260
	13'h0931: q1 = 16'h0c6d; // 0x1262
	13'h0932: q1 = 16'h0049; // 0x1264
	13'h0933: q1 = 16'h0012; // 0x1266
	13'h0934: q1 = 16'h660a; // 0x1268
	13'h0935: q1 = 16'h3b7c; // 0x126a
	13'h0936: q1 = 16'h0001; // 0x126c
	13'h0937: q1 = 16'h0018; // 0x126e
	13'h0938: q1 = 16'h6000; // 0x1270
	13'h0939: q1 = 16'h0220; // 0x1272
	13'h093a: q1 = 16'h0c6d; // 0x1274
	13'h093b: q1 = 16'h000b; // 0x1276
	13'h093c: q1 = 16'h0012; // 0x1278
	13'h093d: q1 = 16'h6e00; // 0x127a
	13'h093e: q1 = 16'h0082; // 0x127c
	13'h093f: q1 = 16'h3a2d; // 0x127e
	13'h0940: q1 = 16'h0012; // 0x1280
	13'h0941: q1 = 16'h5345; // 0x1282
	13'h0942: q1 = 16'h206d; // 0x1284
	13'h0943: q1 = 16'h0024; // 0x1286
	13'h0944: q1 = 16'h3205; // 0x1288
	13'h0945: q1 = 16'h48c1; // 0x128a
	13'h0946: q1 = 16'hd2bc; // 0x128c
	13'h0947: q1 = 16'h0000; // 0x128e
	13'h0948: q1 = 16'hcb22; // 0x1290
	13'h0949: q1 = 16'h2241; // 0x1292
	13'h094a: q1 = 16'h1211; // 0x1294
	13'h094b: q1 = 16'h4881; // 0x1296
	13'h094c: q1 = 16'h3141; // 0x1298
	13'h094d: q1 = 16'h0004; // 0x129a
	13'h094e: q1 = 16'h206d; // 0x129c
	13'h094f: q1 = 16'h0020; // 0x129e
	13'h0950: q1 = 16'h3205; // 0x12a0
	13'h0951: q1 = 16'h48c1; // 0x12a2
	13'h0952: q1 = 16'hd2bc; // 0x12a4
	13'h0953: q1 = 16'h0000; // 0x12a6
	13'h0954: q1 = 16'hcb2e; // 0x12a8
	13'h0955: q1 = 16'h2241; // 0x12aa
	13'h0956: q1 = 16'h1211; // 0x12ac
	13'h0957: q1 = 16'h4881; // 0x12ae
	13'h0958: q1 = 16'h3141; // 0x12b0
	13'h0959: q1 = 16'h0004; // 0x12b2
	13'h095a: q1 = 16'h206d; // 0x12b4
	13'h095b: q1 = 16'h002c; // 0x12b6
	13'h095c: q1 = 16'h3205; // 0x12b8
	13'h095d: q1 = 16'h48c1; // 0x12ba
	13'h095e: q1 = 16'hd2bc; // 0x12bc
	13'h095f: q1 = 16'h0000; // 0x12be
	13'h0960: q1 = 16'hcb3a; // 0x12c0
	13'h0961: q1 = 16'h2241; // 0x12c2
	13'h0962: q1 = 16'h1211; // 0x12c4
	13'h0963: q1 = 16'h4881; // 0x12c6
	13'h0964: q1 = 16'h3141; // 0x12c8
	13'h0965: q1 = 16'h0004; // 0x12ca
	13'h0966: q1 = 16'h206d; // 0x12cc
	13'h0967: q1 = 16'h0028; // 0x12ce
	13'h0968: q1 = 16'h3205; // 0x12d0
	13'h0969: q1 = 16'h48c1; // 0x12d2
	13'h096a: q1 = 16'hd2bc; // 0x12d4
	13'h096b: q1 = 16'h0000; // 0x12d6
	13'h096c: q1 = 16'hcb46; // 0x12d8
	13'h096d: q1 = 16'h2241; // 0x12da
	13'h096e: q1 = 16'h1211; // 0x12dc
	13'h096f: q1 = 16'h4881; // 0x12de
	13'h0970: q1 = 16'h3141; // 0x12e0
	13'h0971: q1 = 16'h0004; // 0x12e2
	13'h0972: q1 = 16'h303c; // 0x12e4
	13'h0973: q1 = 16'h0100; // 0x12e6
	13'h0974: q1 = 16'h226d; // 0x12e8
	13'h0975: q1 = 16'h0020; // 0x12ea
	13'h0976: q1 = 16'h9169; // 0x12ec
	13'h0977: q1 = 16'h0002; // 0x12ee
	13'h0978: q1 = 16'h206d; // 0x12f0
	13'h0979: q1 = 16'h002c; // 0x12f2
	13'h097a: q1 = 16'h226d; // 0x12f4
	13'h097b: q1 = 16'h0020; // 0x12f6
	13'h097c: q1 = 16'h3169; // 0x12f8
	13'h097d: q1 = 16'h0002; // 0x12fa
	13'h097e: q1 = 16'h0002; // 0x12fc
	13'h097f: q1 = 16'h0c6d; // 0x12fe
	13'h0980: q1 = 16'h0001; // 0x1300
	13'h0981: q1 = 16'h0012; // 0x1302
	13'h0982: q1 = 16'h660c; // 0x1304
	13'h0983: q1 = 16'h2ebc; // 0x1306
	13'h0984: q1 = 16'h0000; // 0x1308
	13'h0985: q1 = 16'hc972; // 0x130a
	13'h0986: q1 = 16'h4eb9; // 0x130c
	13'h0987: q1 = 16'h0000; // 0x130e
	13'h0988: q1 = 16'h7dd8; // 0x1310
	13'h0989: q1 = 16'h0c6d; // 0x1312
	13'h098a: q1 = 16'h0023; // 0x1314
	13'h098b: q1 = 16'h0012; // 0x1316
	13'h098c: q1 = 16'h6628; // 0x1318
	13'h098d: q1 = 16'h2079; // 0x131a
	13'h098e: q1 = 16'h0001; // 0x131c
	13'h098f: q1 = 16'h7fb8; // 0x131e
	13'h0990: q1 = 16'h0c68; // 0x1320
	13'h0991: q1 = 16'h0001; // 0x1322
	13'h0992: q1 = 16'h0002; // 0x1324
	13'h0993: q1 = 16'h660e; // 0x1326
	13'h0994: q1 = 16'h2ebc; // 0x1328
	13'h0995: q1 = 16'h0000; // 0x132a
	13'h0996: q1 = 16'hc674; // 0x132c
	13'h0997: q1 = 16'h4eb9; // 0x132e
	13'h0998: q1 = 16'h0000; // 0x1330
	13'h0999: q1 = 16'h7ff8; // 0x1332
	13'h099a: q1 = 16'h600c; // 0x1334
	13'h099b: q1 = 16'h2ebc; // 0x1336
	13'h099c: q1 = 16'h0000; // 0x1338
	13'h099d: q1 = 16'hc6f2; // 0x133a
	13'h099e: q1 = 16'h4eb9; // 0x133c
	13'h099f: q1 = 16'h0000; // 0x133e
	13'h09a0: q1 = 16'h7ff8; // 0x1340
	13'h09a1: q1 = 16'h526d; // 0x1342
	13'h09a2: q1 = 16'h0012; // 0x1344
	13'h09a3: q1 = 16'h0c6d; // 0x1346
	13'h09a4: q1 = 16'h0002; // 0x1348
	13'h09a5: q1 = 16'h001a; // 0x134a
	13'h09a6: q1 = 16'h6600; // 0x134c
	13'h09a7: q1 = 16'h008a; // 0x134e
	13'h09a8: q1 = 16'h0c6d; // 0x1350
	13'h09a9: q1 = 16'h0025; // 0x1352
	13'h09aa: q1 = 16'h0012; // 0x1354
	13'h09ab: q1 = 16'h661e; // 0x1356
	13'h09ac: q1 = 16'h3b7c; // 0x1358
	13'h09ad: q1 = 16'h0001; // 0x135a
	13'h09ae: q1 = 16'h0018; // 0x135c
	13'h09af: q1 = 16'h206d; // 0x135e
	13'h09b0: q1 = 16'h0020; // 0x1360
	13'h09b1: q1 = 16'h317c; // 0x1362
	13'h09b2: q1 = 16'h008c; // 0x1364
	13'h09b3: q1 = 16'h0004; // 0x1366
	13'h09b4: q1 = 16'h206d; // 0x1368
	13'h09b5: q1 = 16'h002c; // 0x136a
	13'h09b6: q1 = 16'h317c; // 0x136c
	13'h09b7: q1 = 16'h00cc; // 0x136e
	13'h09b8: q1 = 16'h0004; // 0x1370
	13'h09b9: q1 = 16'h6000; // 0x1372
	13'h09ba: q1 = 16'h011e; // 0x1374
	13'h09bb: q1 = 16'h506d; // 0x1376
	13'h09bc: q1 = 16'h000e; // 0x1378
	13'h09bd: q1 = 16'h0c6d; // 0x137a
	13'h09be: q1 = 16'h0047; // 0x137c
	13'h09bf: q1 = 16'h000e; // 0x137e
	13'h09c0: q1 = 16'h6f06; // 0x1380
	13'h09c1: q1 = 16'h046d; // 0x1382
	13'h09c2: q1 = 16'h0048; // 0x1384
	13'h09c3: q1 = 16'h000e; // 0x1386
	13'h09c4: q1 = 16'h206d; // 0x1388
	13'h09c5: q1 = 16'h0024; // 0x138a
	13'h09c6: q1 = 16'h317c; // 0x138c
	13'h09c7: q1 = 16'h00bf; // 0x138e
	13'h09c8: q1 = 16'h0004; // 0x1390
	13'h09c9: q1 = 16'h206d; // 0x1392
	13'h09ca: q1 = 16'h0028; // 0x1394
	13'h09cb: q1 = 16'h317c; // 0x1396
	13'h09cc: q1 = 16'h00be; // 0x1398
	13'h09cd: q1 = 16'h0004; // 0x139a
	13'h09ce: q1 = 16'h302d; // 0x139c
	13'h09cf: q1 = 16'h000e; // 0x139e
	13'h09d0: q1 = 16'h48c0; // 0x13a0
	13'h09d1: q1 = 16'hd0bc; // 0x13a2
	13'h09d2: q1 = 16'h0000; // 0x13a4
	13'h09d3: q1 = 16'hca18; // 0x13a6
	13'h09d4: q1 = 16'h2040; // 0x13a8
	13'h09d5: q1 = 16'h1e10; // 0x13aa
	13'h09d6: q1 = 16'h4887; // 0x13ac
	13'h09d7: q1 = 16'h206d; // 0x13ae
	13'h09d8: q1 = 16'h0020; // 0x13b0
	13'h09d9: q1 = 16'h3207; // 0x13b2
	13'h09da: q1 = 16'hd27c; // 0x13b4
	13'h09db: q1 = 16'h000c; // 0x13b6
	13'h09dc: q1 = 16'h3141; // 0x13b8
	13'h09dd: q1 = 16'h0004; // 0x13ba
	13'h09de: q1 = 16'h206d; // 0x13bc
	13'h09df: q1 = 16'h002c; // 0x13be
	13'h09e0: q1 = 16'h3207; // 0x13c0
	13'h09e1: q1 = 16'h48c1; // 0x13c2
	13'h09e2: q1 = 16'hd2bc; // 0x13c4
	13'h09e3: q1 = 16'h0000; // 0x13c6
	13'h09e4: q1 = 16'hcb62; // 0x13c8
	13'h09e5: q1 = 16'h2241; // 0x13ca
	13'h09e6: q1 = 16'h1211; // 0x13cc
	13'h09e7: q1 = 16'h4881; // 0x13ce
	13'h09e8: q1 = 16'h3141; // 0x13d0
	13'h09e9: q1 = 16'h0004; // 0x13d2
	13'h09ea: q1 = 16'h526d; // 0x13d4
	13'h09eb: q1 = 16'h0012; // 0x13d6
	13'h09ec: q1 = 16'h0c6d; // 0x13d8
	13'h09ed: q1 = 16'h0003; // 0x13da
	13'h09ee: q1 = 16'h001a; // 0x13dc
	13'h09ef: q1 = 16'h6616; // 0x13de
	13'h09f0: q1 = 16'h0c6d; // 0x13e0
	13'h09f1: q1 = 16'h0025; // 0x13e2
	13'h09f2: q1 = 16'h0012; // 0x13e4
	13'h09f3: q1 = 16'h660a; // 0x13e6
	13'h09f4: q1 = 16'h3b7c; // 0x13e8
	13'h09f5: q1 = 16'h0001; // 0x13ea
	13'h09f6: q1 = 16'h0018; // 0x13ec
	13'h09f7: q1 = 16'h6000; // 0x13ee
	13'h09f8: q1 = 16'h00a2; // 0x13f0
	13'h09f9: q1 = 16'h526d; // 0x13f2
	13'h09fa: q1 = 16'h0012; // 0x13f4
	13'h09fb: q1 = 16'h0c6d; // 0x13f6
	13'h09fc: q1 = 16'h0004; // 0x13f8
	13'h09fd: q1 = 16'h001a; // 0x13fa
	13'h09fe: q1 = 16'h6600; // 0x13fc
	13'h09ff: q1 = 16'h0094; // 0x13fe
	13'h0a00: q1 = 16'h206d; // 0x1400
	13'h0a01: q1 = 16'h0024; // 0x1402
	13'h0a02: q1 = 16'h3e10; // 0x1404
	13'h0a03: q1 = 16'hde7c; // 0x1406
	13'h0a04: q1 = 16'hc380; // 0x1408
	13'h0a05: q1 = 16'h4a47; // 0x140a
	13'h0a06: q1 = 16'h6c06; // 0x140c
	13'h0a07: q1 = 16'h3007; // 0x140e
	13'h0a08: q1 = 16'h4440; // 0x1410
	13'h0a09: q1 = 16'h3e00; // 0x1412
	13'h0a0a: q1 = 16'h206d; // 0x1414
	13'h0a0b: q1 = 16'h0024; // 0x1416
	13'h0a0c: q1 = 16'h3c28; // 0x1418
	13'h0a0d: q1 = 16'h0002; // 0x141a
	13'h0a0e: q1 = 16'hdc7c; // 0x141c
	13'h0a0f: q1 = 16'hbc00; // 0x141e
	13'h0a10: q1 = 16'h4a46; // 0x1420
	13'h0a11: q1 = 16'h6c06; // 0x1422
	13'h0a12: q1 = 16'h3006; // 0x1424
	13'h0a13: q1 = 16'h4440; // 0x1426
	13'h0a14: q1 = 16'h3c00; // 0x1428
	13'h0a15: q1 = 16'hbe7c; // 0x142a
	13'h0a16: q1 = 16'h0400; // 0x142c
	13'h0a17: q1 = 16'h6c06; // 0x142e
	13'h0a18: q1 = 16'hbc7c; // 0x1430
	13'h0a19: q1 = 16'h0400; // 0x1432
	13'h0a1a: q1 = 16'h6d06; // 0x1434
	13'h0a1b: q1 = 16'h4a6d; // 0x1436
	13'h0a1c: q1 = 16'h0010; // 0x1438
	13'h0a1d: q1 = 16'h6630; // 0x143a
	13'h0a1e: q1 = 16'h206d; // 0x143c
	13'h0a1f: q1 = 16'h0020; // 0x143e
	13'h0a20: q1 = 16'h317c; // 0x1440
	13'h0a21: q1 = 16'h008c; // 0x1442
	13'h0a22: q1 = 16'h0004; // 0x1444
	13'h0a23: q1 = 16'h206d; // 0x1446
	13'h0a24: q1 = 16'h002c; // 0x1448
	13'h0a25: q1 = 16'h317c; // 0x144a
	13'h0a26: q1 = 16'h00cc; // 0x144c
	13'h0a27: q1 = 16'h0004; // 0x144e
	13'h0a28: q1 = 16'h206d; // 0x1450
	13'h0a29: q1 = 16'h0024; // 0x1452
	13'h0a2a: q1 = 16'h317c; // 0x1454
	13'h0a2b: q1 = 16'h00bf; // 0x1456
	13'h0a2c: q1 = 16'h0004; // 0x1458
	13'h0a2d: q1 = 16'h206d; // 0x145a
	13'h0a2e: q1 = 16'h0028; // 0x145c
	13'h0a2f: q1 = 16'h317c; // 0x145e
	13'h0a30: q1 = 16'h00be; // 0x1460
	13'h0a31: q1 = 16'h0004; // 0x1462
	13'h0a32: q1 = 16'h3b7c; // 0x1464
	13'h0a33: q1 = 16'h0001; // 0x1466
	13'h0a34: q1 = 16'h0018; // 0x1468
	13'h0a35: q1 = 16'h6026; // 0x146a
	13'h0a36: q1 = 16'h3ebc; // 0x146c
	13'h0a37: q1 = 16'h4400; // 0x146e
	13'h0a38: q1 = 16'h206d; // 0x1470
	13'h0a39: q1 = 16'h0024; // 0x1472
	13'h0a3a: q1 = 16'h3028; // 0x1474
	13'h0a3b: q1 = 16'h0002; // 0x1476
	13'h0a3c: q1 = 16'h9157; // 0x1478
	13'h0a3d: q1 = 16'h3f3c; // 0x147a
	13'h0a3e: q1 = 16'h3c80; // 0x147c
	13'h0a3f: q1 = 16'h206d; // 0x147e
	13'h0a40: q1 = 16'h0024; // 0x1480
	13'h0a41: q1 = 16'h3010; // 0x1482
	13'h0a42: q1 = 16'h9157; // 0x1484
	13'h0a43: q1 = 16'h4eb9; // 0x1486
	13'h0a44: q1 = 16'h0000; // 0x1488
	13'h0a45: q1 = 16'h0a1c; // 0x148a
	13'h0a46: q1 = 16'h4a5f; // 0x148c
	13'h0a47: q1 = 16'h3b40; // 0x148e
	13'h0a48: q1 = 16'h000e; // 0x1490
	13'h0a49: q1 = 16'h4a9f; // 0x1492
	13'h0a4a: q1 = 16'h4cdf; // 0x1494
	13'h0a4b: q1 = 16'h20e0; // 0x1496
	13'h0a4c: q1 = 16'h4e5e; // 0x1498
	13'h0a4d: q1 = 16'h4e75; // 0x149a
	13'h0a4e: q1 = 16'h4e56; // 0x149c
	13'h0a4f: q1 = 16'hffde; // 0x149e
	13'h0a50: q1 = 16'h48e7; // 0x14a0
	13'h0a51: q1 = 16'h1f00; // 0x14a2
	13'h0a52: q1 = 16'h4244; // 0x14a4
	13'h0a53: q1 = 16'h2079; // 0x14a6
	13'h0a54: q1 = 16'h0001; // 0x14a8
	13'h0a55: q1 = 16'h7fb8; // 0x14aa
	13'h0a56: q1 = 16'h3a28; // 0x14ac
	13'h0a57: q1 = 16'h0002; // 0x14ae
	13'h0a58: q1 = 16'h5345; // 0x14b0
	13'h0a59: q1 = 16'hba6e; // 0x14b2
	13'h0a5a: q1 = 16'h0008; // 0x14b4
	13'h0a5b: q1 = 16'h6f40; // 0x14b6
	13'h0a5c: q1 = 16'h200e; // 0x14b8
	13'h0a5d: q1 = 16'hd0bc; // 0x14ba
	13'h0a5e: q1 = 16'hffff; // 0x14bc
	13'h0a5f: q1 = 16'hffe0; // 0x14be
	13'h0a60: q1 = 16'h2e80; // 0x14c0
	13'h0a61: q1 = 16'h3f05; // 0x14c2
	13'h0a62: q1 = 16'h4eb9; // 0x14c4
	13'h0a63: q1 = 16'h0000; // 0x14c6
	13'h0a64: q1 = 16'h0828; // 0x14c8
	13'h0a65: q1 = 16'h4a5f; // 0x14ca
	13'h0a66: q1 = 16'h2ebc; // 0x14cc
	13'h0a67: q1 = 16'h0000; // 0x14ce
	13'h0a68: q1 = 16'hcb20; // 0x14d0
	13'h0a69: q1 = 16'h200e; // 0x14d2
	13'h0a6a: q1 = 16'hd0bc; // 0x14d4
	13'h0a6b: q1 = 16'hffff; // 0x14d6
	13'h0a6c: q1 = 16'hffe0; // 0x14d8
	13'h0a6d: q1 = 16'h2f00; // 0x14da
	13'h0a6e: q1 = 16'h4eb9; // 0x14dc
	13'h0a6f: q1 = 16'h0000; // 0x14de
	13'h0a70: q1 = 16'h0770; // 0x14e0
	13'h0a71: q1 = 16'h4a9f; // 0x14e2
	13'h0a72: q1 = 16'h200e; // 0x14e4
	13'h0a73: q1 = 16'hd0bc; // 0x14e6
	13'h0a74: q1 = 16'hffff; // 0x14e8
	13'h0a75: q1 = 16'hffe0; // 0x14ea
	13'h0a76: q1 = 16'h2e80; // 0x14ec
	13'h0a77: q1 = 16'h4eb9; // 0x14ee
	13'h0a78: q1 = 16'h0000; // 0x14f0
	13'h0a79: q1 = 16'h072e; // 0x14f2
	13'h0a7a: q1 = 16'h3800; // 0x14f4
	13'h0a7b: q1 = 16'h7a01; // 0x14f6
	13'h0a7c: q1 = 16'h4247; // 0x14f8
	13'h0a7d: q1 = 16'hbe45; // 0x14fa
	13'h0a7e: q1 = 16'h6c24; // 0x14fc
	13'h0a7f: q1 = 16'h3004; // 0x14fe
	13'h0a80: q1 = 16'h48c0; // 0x1500
	13'h0a81: q1 = 16'hd08e; // 0x1502
	13'h0a82: q1 = 16'h2040; // 0x1504
	13'h0a83: q1 = 16'h117c; // 0x1506
	13'h0a84: q1 = 16'h0014; // 0x1508
	13'h0a85: q1 = 16'hffe0; // 0x150a
	13'h0a86: q1 = 16'h5244; // 0x150c
	13'h0a87: q1 = 16'h3004; // 0x150e
	13'h0a88: q1 = 16'h48c0; // 0x1510
	13'h0a89: q1 = 16'hd08e; // 0x1512
	13'h0a8a: q1 = 16'h2040; // 0x1514
	13'h0a8b: q1 = 16'h117c; // 0x1516
	13'h0a8c: q1 = 16'h0015; // 0x1518
	13'h0a8d: q1 = 16'hffe0; // 0x151a
	13'h0a8e: q1 = 16'h5244; // 0x151c
	13'h0a8f: q1 = 16'h5247; // 0x151e
	13'h0a90: q1 = 16'h60d8; // 0x1520
	13'h0a91: q1 = 16'h4247; // 0x1522
	13'h0a92: q1 = 16'h302e; // 0x1524
	13'h0a93: q1 = 16'h0008; // 0x1526
	13'h0a94: q1 = 16'he340; // 0x1528
	13'h0a95: q1 = 16'h9044; // 0x152a
	13'h0a96: q1 = 16'hb047; // 0x152c
	13'h0a97: q1 = 16'h6f26; // 0x152e
	13'h0a98: q1 = 16'h7020; // 0x1530
	13'h0a99: q1 = 16'h322e; // 0x1532
	13'h0a9a: q1 = 16'h0008; // 0x1534
	13'h0a9b: q1 = 16'he341; // 0x1536
	13'h0a9c: q1 = 16'h9041; // 0x1538
	13'h0a9d: q1 = 16'h3c00; // 0x153a
	13'h0a9e: q1 = 16'hdc47; // 0x153c
	13'h0a9f: q1 = 16'h4257; // 0x153e
	13'h0aa0: q1 = 16'h3f3c; // 0x1540
	13'h0aa1: q1 = 16'h0040; // 0x1542
	13'h0aa2: q1 = 16'h3f3c; // 0x1544
	13'h0aa3: q1 = 16'h0004; // 0x1546
	13'h0aa4: q1 = 16'h3f06; // 0x1548
	13'h0aa5: q1 = 16'h4eb9; // 0x154a
	13'h0aa6: q1 = 16'h0000; // 0x154c
	13'h0aa7: q1 = 16'h3d18; // 0x154e
	13'h0aa8: q1 = 16'h5c4f; // 0x1550
	13'h0aa9: q1 = 16'h5247; // 0x1552
	13'h0aaa: q1 = 16'h60ce; // 0x1554
	13'h0aab: q1 = 16'h4247; // 0x1556
	13'h0aac: q1 = 16'hbe44; // 0x1558
	13'h0aad: q1 = 16'h6c68; // 0x155a
	13'h0aae: q1 = 16'h7c20; // 0x155c
	13'h0aaf: q1 = 16'h9c44; // 0x155e
	13'h0ab0: q1 = 16'hdc47; // 0x1560
	13'h0ab1: q1 = 16'h3207; // 0x1562
	13'h0ab2: q1 = 16'h48c1; // 0x1564
	13'h0ab3: q1 = 16'h200e; // 0x1566
	13'h0ab4: q1 = 16'hd081; // 0x1568
	13'h0ab5: q1 = 16'h2040; // 0x156a
	13'h0ab6: q1 = 16'h0c28; // 0x156c
	13'h0ab7: q1 = 16'h0014; // 0x156e
	13'h0ab8: q1 = 16'hffe0; // 0x1570
	13'h0ab9: q1 = 16'h6608; // 0x1572
	13'h0aba: q1 = 16'h3d7c; // 0x1574
	13'h0abb: q1 = 16'h0007; // 0x1576
	13'h0abc: q1 = 16'hffde; // 0x1578
	13'h0abd: q1 = 16'h6020; // 0x157a
	13'h0abe: q1 = 16'h3207; // 0x157c
	13'h0abf: q1 = 16'h48c1; // 0x157e
	13'h0ac0: q1 = 16'h200e; // 0x1580
	13'h0ac1: q1 = 16'hd081; // 0x1582
	13'h0ac2: q1 = 16'h2040; // 0x1584
	13'h0ac3: q1 = 16'h0c28; // 0x1586
	13'h0ac4: q1 = 16'h0015; // 0x1588
	13'h0ac5: q1 = 16'hffe0; // 0x158a
	13'h0ac6: q1 = 16'h6608; // 0x158c
	13'h0ac7: q1 = 16'h3d7c; // 0x158e
	13'h0ac8: q1 = 16'h002b; // 0x1590
	13'h0ac9: q1 = 16'hffde; // 0x1592
	13'h0aca: q1 = 16'h6006; // 0x1594
	13'h0acb: q1 = 16'h3d7c; // 0x1596
	13'h0acc: q1 = 16'h0028; // 0x1598
	13'h0acd: q1 = 16'hffde; // 0x159a
	13'h0ace: q1 = 16'h3eae; // 0x159c
	13'h0acf: q1 = 16'hffde; // 0x159e
	13'h0ad0: q1 = 16'h3207; // 0x15a0
	13'h0ad1: q1 = 16'h48c1; // 0x15a2
	13'h0ad2: q1 = 16'h200e; // 0x15a4
	13'h0ad3: q1 = 16'hd081; // 0x15a6
	13'h0ad4: q1 = 16'h2040; // 0x15a8
	13'h0ad5: q1 = 16'h1028; // 0x15aa
	13'h0ad6: q1 = 16'hffe0; // 0x15ac
	13'h0ad7: q1 = 16'h4880; // 0x15ae
	13'h0ad8: q1 = 16'h3f00; // 0x15b0
	13'h0ad9: q1 = 16'h3f3c; // 0x15b2
	13'h0ada: q1 = 16'h0004; // 0x15b4
	13'h0adb: q1 = 16'h3f06; // 0x15b6
	13'h0adc: q1 = 16'h4eb9; // 0x15b8
	13'h0add: q1 = 16'h0000; // 0x15ba
	13'h0ade: q1 = 16'h3d18; // 0x15bc
	13'h0adf: q1 = 16'h5c4f; // 0x15be
	13'h0ae0: q1 = 16'h5247; // 0x15c0
	13'h0ae1: q1 = 16'h6094; // 0x15c2
	13'h0ae2: q1 = 16'h4a9f; // 0x15c4
	13'h0ae3: q1 = 16'h4cdf; // 0x15c6
	13'h0ae4: q1 = 16'h00f0; // 0x15c8
	13'h0ae5: q1 = 16'h4e5e; // 0x15ca
	13'h0ae6: q1 = 16'h4e75; // 0x15cc
	13'h0ae7: q1 = 16'h4e56; // 0x15ce
	13'h0ae8: q1 = 16'h0000; // 0x15d0
	13'h0ae9: q1 = 16'h48e7; // 0x15d2
	13'h0aea: q1 = 16'h0700; // 0x15d4
	13'h0aeb: q1 = 16'h3e2e; // 0x15d6
	13'h0aec: q1 = 16'h0008; // 0x15d8
	13'h0aed: q1 = 16'h3007; // 0x15da
	13'h0aee: q1 = 16'hc1fc; // 0x15dc
	13'h0aef: q1 = 16'h0003; // 0x15de
	13'h0af0: q1 = 16'h3c00; // 0x15e0
	13'h0af1: q1 = 16'hbc7c; // 0x15e2
	13'h0af2: q1 = 16'h002d; // 0x15e4
	13'h0af3: q1 = 16'h6c1e; // 0x15e6
	13'h0af4: q1 = 16'h3006; // 0x15e8
	13'h0af5: q1 = 16'h48c0; // 0x15ea
	13'h0af6: q1 = 16'hd0bc; // 0x15ec
	13'h0af7: q1 = 16'h0001; // 0x15ee
	13'h0af8: q1 = 16'h7ba8; // 0x15f0
	13'h0af9: q1 = 16'h2040; // 0x15f2
	13'h0afa: q1 = 16'h3206; // 0x15f4
	13'h0afb: q1 = 16'h48c1; // 0x15f6
	13'h0afc: q1 = 16'hd2bc; // 0x15f8
	13'h0afd: q1 = 16'h0000; // 0x15fa
	13'h0afe: q1 = 16'hf8f0; // 0x15fc
	13'h0aff: q1 = 16'h2241; // 0x15fe
	13'h0b00: q1 = 16'h1091; // 0x1600
	13'h0b01: q1 = 16'h5246; // 0x1602
	13'h0b02: q1 = 16'h60dc; // 0x1604
	13'h0b03: q1 = 16'h3c07; // 0x1606
	13'h0b04: q1 = 16'hbc7c; // 0x1608
	13'h0b05: q1 = 16'h000f; // 0x160a
	13'h0b06: q1 = 16'h6c48; // 0x160c
	13'h0b07: q1 = 16'h3006; // 0x160e
	13'h0b08: q1 = 16'he340; // 0x1610
	13'h0b09: q1 = 16'h48c0; // 0x1612
	13'h0b0a: q1 = 16'hd0bc; // 0x1614
	13'h0b0b: q1 = 16'h0001; // 0x1616
	13'h0b0c: q1 = 16'h7efe; // 0x1618
	13'h0b0d: q1 = 16'h2040; // 0x161a
	13'h0b0e: q1 = 16'h3206; // 0x161c
	13'h0b0f: q1 = 16'h48c1; // 0x161e
	13'h0b10: q1 = 16'hd2bc; // 0x1620
	13'h0b11: q1 = 16'h0000; // 0x1622
	13'h0b12: q1 = 16'hf93c; // 0x1624
	13'h0b13: q1 = 16'h2241; // 0x1626
	13'h0b14: q1 = 16'h1211; // 0x1628
	13'h0b15: q1 = 16'h4881; // 0x162a
	13'h0b16: q1 = 16'h3081; // 0x162c
	13'h0b17: q1 = 16'h3006; // 0x162e
	13'h0b18: q1 = 16'he340; // 0x1630
	13'h0b19: q1 = 16'h48c0; // 0x1632
	13'h0b1a: q1 = 16'hd0bc; // 0x1634
	13'h0b1b: q1 = 16'h0000; // 0x1636
	13'h0b1c: q1 = 16'hf91e; // 0x1638
	13'h0b1d: q1 = 16'h2040; // 0x163a
	13'h0b1e: q1 = 16'h3f10; // 0x163c
	13'h0b1f: q1 = 16'h3006; // 0x163e
	13'h0b20: q1 = 16'he540; // 0x1640
	13'h0b21: q1 = 16'h48c0; // 0x1642
	13'h0b22: q1 = 16'hd0bc; // 0x1644
	13'h0b23: q1 = 16'h0001; // 0x1646
	13'h0b24: q1 = 16'h7f64; // 0x1648
	13'h0b25: q1 = 16'h2040; // 0x164a
	13'h0b26: q1 = 16'h301f; // 0x164c
	13'h0b27: q1 = 16'h48c0; // 0x164e
	13'h0b28: q1 = 16'h2080; // 0x1650
	13'h0b29: q1 = 16'h5246; // 0x1652
	13'h0b2a: q1 = 16'h60b2; // 0x1654
	13'h0b2b: q1 = 16'h2ebc; // 0x1656
	13'h0b2c: q1 = 16'h0001; // 0x1658
	13'h0b2d: q1 = 16'h860e; // 0x165a
	13'h0b2e: q1 = 16'h2f39; // 0x165c
	13'h0b2f: q1 = 16'h0001; // 0x165e
	13'h0b30: q1 = 16'h7f64; // 0x1660
	13'h0b31: q1 = 16'h4eb9; // 0x1662
	13'h0b32: q1 = 16'h0000; // 0x1664
	13'h0b33: q1 = 16'h0892; // 0x1666
	13'h0b34: q1 = 16'h4a9f; // 0x1668
	13'h0b35: q1 = 16'h2ebc; // 0x166a
	13'h0b36: q1 = 16'h0000; // 0x166c
	13'h0b37: q1 = 16'hcb70; // 0x166e
	13'h0b38: q1 = 16'h2f3c; // 0x1670
	13'h0b39: q1 = 16'h0001; // 0x1672
	13'h0b3a: q1 = 16'h860e; // 0x1674
	13'h0b3b: q1 = 16'h4eb9; // 0x1676
	13'h0b3c: q1 = 16'h0000; // 0x1678
	13'h0b3d: q1 = 16'h0770; // 0x167a
	13'h0b3e: q1 = 16'h4a9f; // 0x167c
	13'h0b3f: q1 = 16'h4a9f; // 0x167e
	13'h0b40: q1 = 16'h4cdf; // 0x1680
	13'h0b41: q1 = 16'h00c0; // 0x1682
	13'h0b42: q1 = 16'h4e5e; // 0x1684
	13'h0b43: q1 = 16'h4e75; // 0x1686
	13'h0b44: q1 = 16'h4e56; // 0x1688
	13'h0b45: q1 = 16'hfffc; // 0x168a
	13'h0b46: q1 = 16'h48e7; // 0x168c
	13'h0b47: q1 = 16'h071c; // 0x168e
	13'h0b48: q1 = 16'h2a7c; // 0x1690
	13'h0b49: q1 = 16'h0001; // 0x1692
	13'h0b4a: q1 = 16'h7f2c; // 0x1694
	13'h0b4b: q1 = 16'h287c; // 0x1696
	13'h0b4c: q1 = 16'h0001; // 0x1698
	13'h0b4d: q1 = 16'h807a; // 0x169a
	13'h0b4e: q1 = 16'h267c; // 0x169c
	13'h0b4f: q1 = 16'h0001; // 0x169e
	13'h0b50: q1 = 16'h80aa; // 0x16a0
	13'h0b51: q1 = 16'h2d7c; // 0x16a2
	13'h0b52: q1 = 16'h0001; // 0x16a4
	13'h0b53: q1 = 16'h80a2; // 0x16a6
	13'h0b54: q1 = 16'hfffc; // 0x16a8
	13'h0b55: q1 = 16'h0c55; // 0x16aa
	13'h0b56: q1 = 16'h0017; // 0x16ac
	13'h0b57: q1 = 16'h6600; // 0x16ae
	13'h0b58: q1 = 16'h00f0; // 0x16b0
	13'h0b59: q1 = 16'h206d; // 0x16b2
	13'h0b5a: q1 = 16'h0020; // 0x16b4
	13'h0b5b: q1 = 16'h317c; // 0x16b6
	13'h0b5c: q1 = 16'h00d2; // 0x16b8
	13'h0b5d: q1 = 16'h0004; // 0x16ba
	13'h0b5e: q1 = 16'h206d; // 0x16bc
	13'h0b5f: q1 = 16'h0020; // 0x16be
	13'h0b60: q1 = 16'h317c; // 0x16c0
	13'h0b61: q1 = 16'h0007; // 0x16c2
	13'h0b62: q1 = 16'h0006; // 0x16c4
	13'h0b63: q1 = 16'h3ebc; // 0x16c6
	13'h0b64: q1 = 16'h0024; // 0x16c8
	13'h0b65: q1 = 16'h202d; // 0x16ca
	13'h0b66: q1 = 16'h0020; // 0x16cc
	13'h0b67: q1 = 16'h5c80; // 0x16ce
	13'h0b68: q1 = 16'h2f00; // 0x16d0
	13'h0b69: q1 = 16'h4eb9; // 0x16d2
	13'h0b6a: q1 = 16'h0000; // 0x16d4
	13'h0b6b: q1 = 16'h3ee6; // 0x16d6
	13'h0b6c: q1 = 16'h4a9f; // 0x16d8
	13'h0b6d: q1 = 16'h206d; // 0x16da
	13'h0b6e: q1 = 16'h002c; // 0x16dc
	13'h0b6f: q1 = 16'h317c; // 0x16de
	13'h0b70: q1 = 16'h00d5; // 0x16e0
	13'h0b71: q1 = 16'h0004; // 0x16e2
	13'h0b72: q1 = 16'h206d; // 0x16e4
	13'h0b73: q1 = 16'h002c; // 0x16e6
	13'h0b74: q1 = 16'h317c; // 0x16e8
	13'h0b75: q1 = 16'h001d; // 0x16ea
	13'h0b76: q1 = 16'h0006; // 0x16ec
	13'h0b77: q1 = 16'h3ebc; // 0x16ee
	13'h0b78: q1 = 16'h0024; // 0x16f0
	13'h0b79: q1 = 16'h202d; // 0x16f2
	13'h0b7a: q1 = 16'h002c; // 0x16f4
	13'h0b7b: q1 = 16'h5c80; // 0x16f6
	13'h0b7c: q1 = 16'h2f00; // 0x16f8
	13'h0b7d: q1 = 16'h4eb9; // 0x16fa
	13'h0b7e: q1 = 16'h0000; // 0x16fc
	13'h0b7f: q1 = 16'h3ee6; // 0x16fe
	13'h0b80: q1 = 16'h4a9f; // 0x1700
	13'h0b81: q1 = 16'h206d; // 0x1702
	13'h0b82: q1 = 16'h0024; // 0x1704
	13'h0b83: q1 = 16'h3239; // 0x1706
	13'h0b84: q1 = 16'h0001; // 0x1708
	13'h0b85: q1 = 16'h8938; // 0x170a
	13'h0b86: q1 = 16'hd27c; // 0x170c
	13'h0b87: q1 = 16'hfd00; // 0x170e
	13'h0b88: q1 = 16'h3141; // 0x1710
	13'h0b89: q1 = 16'h0002; // 0x1712
	13'h0b8a: q1 = 16'h206d; // 0x1714
	13'h0b8b: q1 = 16'h0024; // 0x1716
	13'h0b8c: q1 = 16'h3b68; // 0x1718
	13'h0b8d: q1 = 16'h0002; // 0x171a
	13'h0b8e: q1 = 16'h0030; // 0x171c
	13'h0b8f: q1 = 16'h206d; // 0x171e
	13'h0b90: q1 = 16'h0020; // 0x1720
	13'h0b91: q1 = 16'h226d; // 0x1722
	13'h0b92: q1 = 16'h0024; // 0x1724
	13'h0b93: q1 = 16'h3091; // 0x1726
	13'h0b94: q1 = 16'h206d; // 0x1728
	13'h0b95: q1 = 16'h0020; // 0x172a
	13'h0b96: q1 = 16'h226d; // 0x172c
	13'h0b97: q1 = 16'h0024; // 0x172e
	13'h0b98: q1 = 16'h3229; // 0x1730
	13'h0b99: q1 = 16'h0002; // 0x1732
	13'h0b9a: q1 = 16'hd27c; // 0x1734
	13'h0b9b: q1 = 16'h0200; // 0x1736
	13'h0b9c: q1 = 16'h3141; // 0x1738
	13'h0b9d: q1 = 16'h0002; // 0x173a
	13'h0b9e: q1 = 16'h206d; // 0x173c
	13'h0b9f: q1 = 16'h002c; // 0x173e
	13'h0ba0: q1 = 16'h226d; // 0x1740
	13'h0ba1: q1 = 16'h0020; // 0x1742
	13'h0ba2: q1 = 16'h3091; // 0x1744
	13'h0ba3: q1 = 16'h206d; // 0x1746
	13'h0ba4: q1 = 16'h002c; // 0x1748
	13'h0ba5: q1 = 16'h226d; // 0x174a
	13'h0ba6: q1 = 16'h0020; // 0x174c
	13'h0ba7: q1 = 16'h3169; // 0x174e
	13'h0ba8: q1 = 16'h0002; // 0x1750
	13'h0ba9: q1 = 16'h0002; // 0x1752
	13'h0baa: q1 = 16'h206d; // 0x1754
	13'h0bab: q1 = 16'h0024; // 0x1756
	13'h0bac: q1 = 16'h317c; // 0x1758
	13'h0bad: q1 = 16'h00bf; // 0x175a
	13'h0bae: q1 = 16'h0004; // 0x175c
	13'h0baf: q1 = 16'h4aad; // 0x175e
	13'h0bb0: q1 = 16'h0006; // 0x1760
	13'h0bb1: q1 = 16'h670c; // 0x1762
	13'h0bb2: q1 = 16'h206d; // 0x1764
	13'h0bb3: q1 = 16'h0028; // 0x1766
	13'h0bb4: q1 = 16'h317c; // 0x1768
	13'h0bb5: q1 = 16'h00f2; // 0x176a
	13'h0bb6: q1 = 16'h0004; // 0x176c
	13'h0bb7: q1 = 16'h600a; // 0x176e
	13'h0bb8: q1 = 16'h206d; // 0x1770
	13'h0bb9: q1 = 16'h0028; // 0x1772
	13'h0bba: q1 = 16'h317c; // 0x1774
	13'h0bbb: q1 = 16'h00be; // 0x1776
	13'h0bbc: q1 = 16'h0004; // 0x1778
	13'h0bbd: q1 = 16'h206d; // 0x177a
	13'h0bbe: q1 = 16'h0028; // 0x177c
	13'h0bbf: q1 = 16'h226d; // 0x177e
	13'h0bc0: q1 = 16'h0024; // 0x1780
	13'h0bc1: q1 = 16'h3091; // 0x1782
	13'h0bc2: q1 = 16'h206d; // 0x1784
	13'h0bc3: q1 = 16'h0028; // 0x1786
	13'h0bc4: q1 = 16'h226d; // 0x1788
	13'h0bc5: q1 = 16'h0024; // 0x178a
	13'h0bc6: q1 = 16'h3169; // 0x178c
	13'h0bc7: q1 = 16'h0002; // 0x178e
	13'h0bc8: q1 = 16'h0002; // 0x1790
	13'h0bc9: q1 = 16'h5255; // 0x1792
	13'h0bca: q1 = 16'h4eb9; // 0x1794
	13'h0bcb: q1 = 16'h0000; // 0x1796
	13'h0bcc: q1 = 16'h4340; // 0x1798
	13'h0bcd: q1 = 16'h7001; // 0x179a
	13'h0bce: q1 = 16'h6000; // 0x179c
	13'h0bcf: q1 = 16'h02f4; // 0x179e
	13'h0bd0: q1 = 16'h3c15; // 0x17a0
	13'h0bd1: q1 = 16'hbc7c; // 0x17a2
	13'h0bd2: q1 = 16'h0007; // 0x17a4
	13'h0bd3: q1 = 16'h6f04; // 0x17a6
	13'h0bd4: q1 = 16'h5146; // 0x17a8
	13'h0bd5: q1 = 16'h60f6; // 0x17aa
	13'h0bd6: q1 = 16'h206d; // 0x17ac
	13'h0bd7: q1 = 16'h0024; // 0x17ae
	13'h0bd8: q1 = 16'h3206; // 0x17b0
	13'h0bd9: q1 = 16'h48c1; // 0x17b2
	13'h0bda: q1 = 16'hd2bc; // 0x17b4
	13'h0bdb: q1 = 16'h0000; // 0x17b6
	13'h0bdc: q1 = 16'hcb5a; // 0x17b8
	13'h0bdd: q1 = 16'h2241; // 0x17ba
	13'h0bde: q1 = 16'h1211; // 0x17bc
	13'h0bdf: q1 = 16'h4881; // 0x17be
	13'h0be0: q1 = 16'h3141; // 0x17c0
	13'h0be1: q1 = 16'h0004; // 0x17c2
	13'h0be2: q1 = 16'h206d; // 0x17c4
	13'h0be3: q1 = 16'h0024; // 0x17c6
	13'h0be4: q1 = 16'h3215; // 0x17c8
	13'h0be5: q1 = 16'h48c1; // 0x17ca
	13'h0be6: q1 = 16'hd2bc; // 0x17cc
	13'h0be7: q1 = 16'h0000; // 0x17ce
	13'h0be8: q1 = 16'hcbec; // 0x17d0
	13'h0be9: q1 = 16'h2241; // 0x17d2
	13'h0bea: q1 = 16'h1211; // 0x17d4
	13'h0beb: q1 = 16'h4881; // 0x17d6
	13'h0bec: q1 = 16'h5f41; // 0x17d8
	13'h0bed: q1 = 16'hef41; // 0x17da
	13'h0bee: q1 = 16'hd279; // 0x17dc
	13'h0bef: q1 = 16'h0001; // 0x17de
	13'h0bf0: q1 = 16'h8936; // 0x17e0
	13'h0bf1: q1 = 16'h3081; // 0x17e2
	13'h0bf2: q1 = 16'h206d; // 0x17e4
	13'h0bf3: q1 = 16'h0024; // 0x17e6
	13'h0bf4: q1 = 16'h3239; // 0x17e8
	13'h0bf5: q1 = 16'h0001; // 0x17ea
	13'h0bf6: q1 = 16'h8938; // 0x17ec
	13'h0bf7: q1 = 16'hd27c; // 0x17ee
	13'h0bf8: q1 = 16'hfd00; // 0x17f0
	13'h0bf9: q1 = 16'h3415; // 0x17f2
	13'h0bfa: q1 = 16'h48c2; // 0x17f4
	13'h0bfb: q1 = 16'hd4bc; // 0x17f6
	13'h0bfc: q1 = 16'h0000; // 0x17f8
	13'h0bfd: q1 = 16'hcc04; // 0x17fa
	13'h0bfe: q1 = 16'h2442; // 0x17fc
	13'h0bff: q1 = 16'h1412; // 0x17fe
	13'h0c00: q1 = 16'h4882; // 0x1800
	13'h0c01: q1 = 16'hef42; // 0x1802
	13'h0c02: q1 = 16'h9242; // 0x1804
	13'h0c03: q1 = 16'h3141; // 0x1806
	13'h0c04: q1 = 16'h0002; // 0x1808
	13'h0c05: q1 = 16'h206d; // 0x180a
	13'h0c06: q1 = 16'h0024; // 0x180c
	13'h0c07: q1 = 16'h0c68; // 0x180e
	13'h0c08: q1 = 16'h1280; // 0x1810
	13'h0c09: q1 = 16'h0002; // 0x1812
	13'h0c0a: q1 = 16'h6c0a; // 0x1814
	13'h0c0b: q1 = 16'h206d; // 0x1816
	13'h0c0c: q1 = 16'h0024; // 0x1818
	13'h0c0d: q1 = 16'h317c; // 0x181a
	13'h0c0e: q1 = 16'h1280; // 0x181c
	13'h0c0f: q1 = 16'h0002; // 0x181e
	13'h0c10: q1 = 16'h206d; // 0x1820
	13'h0c11: q1 = 16'h0024; // 0x1822
	13'h0c12: q1 = 16'h3b68; // 0x1824
	13'h0c13: q1 = 16'h0002; // 0x1826
	13'h0c14: q1 = 16'h0030; // 0x1828
	13'h0c15: q1 = 16'h4eb9; // 0x182a
	13'h0c16: q1 = 16'h0000; // 0x182c
	13'h0c17: q1 = 16'h607a; // 0x182e
	13'h0c18: q1 = 16'h4aad; // 0x1830
	13'h0c19: q1 = 16'h0006; // 0x1832
	13'h0c1a: q1 = 16'h670c; // 0x1834
	13'h0c1b: q1 = 16'h206d; // 0x1836
	13'h0c1c: q1 = 16'h0028; // 0x1838
	13'h0c1d: q1 = 16'h317c; // 0x183a
	13'h0c1e: q1 = 16'h00f2; // 0x183c
	13'h0c1f: q1 = 16'h0004; // 0x183e
	13'h0c20: q1 = 16'h6018; // 0x1840
	13'h0c21: q1 = 16'h206d; // 0x1842
	13'h0c22: q1 = 16'h0028; // 0x1844
	13'h0c23: q1 = 16'h3206; // 0x1846
	13'h0c24: q1 = 16'h48c1; // 0x1848
	13'h0c25: q1 = 16'hd2bc; // 0x184a
	13'h0c26: q1 = 16'h0000; // 0x184c
	13'h0c27: q1 = 16'hcb52; // 0x184e
	13'h0c28: q1 = 16'h2241; // 0x1850
	13'h0c29: q1 = 16'h1211; // 0x1852
	13'h0c2a: q1 = 16'h4881; // 0x1854
	13'h0c2b: q1 = 16'h3141; // 0x1856
	13'h0c2c: q1 = 16'h0004; // 0x1858
	13'h0c2d: q1 = 16'hbc7c; // 0x185a
	13'h0c2e: q1 = 16'h0001; // 0x185c
	13'h0c2f: q1 = 16'h6706; // 0x185e
	13'h0c30: q1 = 16'hbc7c; // 0x1860
	13'h0c31: q1 = 16'h0005; // 0x1862
	13'h0c32: q1 = 16'h6614; // 0x1864
	13'h0c33: q1 = 16'h4a79; // 0x1866
	13'h0c34: q1 = 16'h0001; // 0x1868
	13'h0c35: q1 = 16'h8676; // 0x186a
	13'h0c36: q1 = 16'h660c; // 0x186c
	13'h0c37: q1 = 16'h2ebc; // 0x186e
	13'h0c38: q1 = 16'h0000; // 0x1870
	13'h0c39: q1 = 16'hfd1c; // 0x1872
	13'h0c3a: q1 = 16'h4eb9; // 0x1874
	13'h0c3b: q1 = 16'h0000; // 0x1876
	13'h0c3c: q1 = 16'h7dd8; // 0x1878
	13'h0c3d: q1 = 16'h3015; // 0x187a
	13'h0c3e: q1 = 16'h48c0; // 0x187c
	13'h0c3f: q1 = 16'hd0bc; // 0x187e
	13'h0c40: q1 = 16'h0000; // 0x1880
	13'h0c41: q1 = 16'hcb74; // 0x1882
	13'h0c42: q1 = 16'h2040; // 0x1884
	13'h0c43: q1 = 16'h1010; // 0x1886
	13'h0c44: q1 = 16'h4880; // 0x1888
	13'h0c45: q1 = 16'h3940; // 0x188a
	13'h0c46: q1 = 16'h0004; // 0x188c
	13'h0c47: q1 = 16'h397c; // 0x188e
	13'h0c48: q1 = 16'h000d; // 0x1890
	13'h0c49: q1 = 16'h0006; // 0x1892
	13'h0c4a: q1 = 16'h206d; // 0x1894
	13'h0c4b: q1 = 16'h0024; // 0x1896
	13'h0c4c: q1 = 16'h3890; // 0x1898
	13'h0c4d: q1 = 16'h206d; // 0x189a
	13'h0c4e: q1 = 16'h0024; // 0x189c
	13'h0c4f: q1 = 16'h3028; // 0x189e
	13'h0c50: q1 = 16'h0002; // 0x18a0
	13'h0c51: q1 = 16'h3215; // 0x18a2
	13'h0c52: q1 = 16'h48c1; // 0x18a4
	13'h0c53: q1 = 16'hd2bc; // 0x18a6
	13'h0c54: q1 = 16'h0000; // 0x18a8
	13'h0c55: q1 = 16'hcc04; // 0x18aa
	13'h0c56: q1 = 16'h2241; // 0x18ac
	13'h0c57: q1 = 16'h1211; // 0x18ae
	13'h0c58: q1 = 16'h4881; // 0x18b0
	13'h0c59: q1 = 16'hef41; // 0x18b2
	13'h0c5a: q1 = 16'hd041; // 0x18b4
	13'h0c5b: q1 = 16'hd07c; // 0x18b6
	13'h0c5c: q1 = 16'h0380; // 0x18b8
	13'h0c5d: q1 = 16'h3940; // 0x18ba
	13'h0c5e: q1 = 16'h0002; // 0x18bc
	13'h0c5f: q1 = 16'h0c55; // 0x18be
	13'h0c60: q1 = 16'h0002; // 0x18c0
	13'h0c61: q1 = 16'h6f00; // 0x18c2
	13'h0c62: q1 = 16'h010c; // 0x18c4
	13'h0c63: q1 = 16'h0c55; // 0x18c6
	13'h0c64: q1 = 16'h0014; // 0x18c8
	13'h0c65: q1 = 16'h6c00; // 0x18ca
	13'h0c66: q1 = 16'h0104; // 0x18cc
	13'h0c67: q1 = 16'h206d; // 0x18ce
	13'h0c68: q1 = 16'h0024; // 0x18d0
	13'h0c69: q1 = 16'h3010; // 0x18d2
	13'h0c6a: q1 = 16'hd07c; // 0x18d4
	13'h0c6b: q1 = 16'hfc00; // 0x18d6
	13'h0c6c: q1 = 16'h3880; // 0x18d8
	13'h0c6d: q1 = 16'h206d; // 0x18da
	13'h0c6e: q1 = 16'h0024; // 0x18dc
	13'h0c6f: q1 = 16'h3028; // 0x18de
	13'h0c70: q1 = 16'h0002; // 0x18e0
	13'h0c71: q1 = 16'h3215; // 0x18e2
	13'h0c72: q1 = 16'h48c1; // 0x18e4
	13'h0c73: q1 = 16'hd2bc; // 0x18e6
	13'h0c74: q1 = 16'h0000; // 0x18e8
	13'h0c75: q1 = 16'hcc04; // 0x18ea
	13'h0c76: q1 = 16'h2241; // 0x18ec
	13'h0c77: q1 = 16'h1211; // 0x18ee
	13'h0c78: q1 = 16'h4881; // 0x18f0
	13'h0c79: q1 = 16'hef41; // 0x18f2
	13'h0c7a: q1 = 16'hd041; // 0x18f4
	13'h0c7b: q1 = 16'hd07c; // 0x18f6
	13'h0c7c: q1 = 16'h0780; // 0x18f8
	13'h0c7d: q1 = 16'h3940; // 0x18fa
	13'h0c7e: q1 = 16'h0002; // 0x18fc
	13'h0c7f: q1 = 16'h396c; // 0x18fe
	13'h0c80: q1 = 16'h0002; // 0x1900
	13'h0c81: q1 = 16'h000a; // 0x1902
	13'h0c82: q1 = 16'h302c; // 0x1904
	13'h0c83: q1 = 16'h0002; // 0x1906
	13'h0c84: q1 = 16'hd07c; // 0x1908
	13'h0c85: q1 = 16'hf800; // 0x190a
	13'h0c86: q1 = 16'h3940; // 0x190c
	13'h0c87: q1 = 16'h0012; // 0x190e
	13'h0c88: q1 = 16'h396c; // 0x1910
	13'h0c89: q1 = 16'h0012; // 0x1912
	13'h0c8a: q1 = 16'h001a; // 0x1914
	13'h0c8b: q1 = 16'h0c55; // 0x1916
	13'h0c8c: q1 = 16'h000b; // 0x1918
	13'h0c8d: q1 = 16'h6f08; // 0x191a
	13'h0c8e: q1 = 16'h376c; // 0x191c
	13'h0c8f: q1 = 16'h0002; // 0x191e
	13'h0c90: q1 = 16'h0002; // 0x1920
	13'h0c91: q1 = 16'h6006; // 0x1922
	13'h0c92: q1 = 16'h376c; // 0x1924
	13'h0c93: q1 = 16'h0012; // 0x1926
	13'h0c94: q1 = 16'h0002; // 0x1928
	13'h0c95: q1 = 16'h3014; // 0x192a
	13'h0c96: q1 = 16'hd07c; // 0x192c
	13'h0c97: q1 = 16'h0800; // 0x192e
	13'h0c98: q1 = 16'h3940; // 0x1930
	13'h0c99: q1 = 16'h0008; // 0x1932
	13'h0c9a: q1 = 16'h3954; // 0x1934
	13'h0c9b: q1 = 16'h0010; // 0x1936
	13'h0c9c: q1 = 16'h396c; // 0x1938
	13'h0c9d: q1 = 16'h0008; // 0x193a
	13'h0c9e: q1 = 16'h0018; // 0x193c
	13'h0c9f: q1 = 16'h0c55; // 0x193e
	13'h0ca0: q1 = 16'h000b; // 0x1940
	13'h0ca1: q1 = 16'h6f04; // 0x1942
	13'h0ca2: q1 = 16'h3694; // 0x1944
	13'h0ca3: q1 = 16'h6008; // 0x1946
	13'h0ca4: q1 = 16'h3014; // 0x1948
	13'h0ca5: q1 = 16'hd07c; // 0x194a
	13'h0ca6: q1 = 16'hf800; // 0x194c
	13'h0ca7: q1 = 16'h3680; // 0x194e
	13'h0ca8: q1 = 16'h3015; // 0x1950
	13'h0ca9: q1 = 16'h48c0; // 0x1952
	13'h0caa: q1 = 16'hd0bc; // 0x1954
	13'h0cab: q1 = 16'h0000; // 0x1956
	13'h0cac: q1 = 16'hcb74; // 0x1958
	13'h0cad: q1 = 16'h2040; // 0x195a
	13'h0cae: q1 = 16'h1010; // 0x195c
	13'h0caf: q1 = 16'h4880; // 0x195e
	13'h0cb0: q1 = 16'h5240; // 0x1960
	13'h0cb1: q1 = 16'h3940; // 0x1962
	13'h0cb2: q1 = 16'h000c; // 0x1964
	13'h0cb3: q1 = 16'h3015; // 0x1966
	13'h0cb4: q1 = 16'h48c0; // 0x1968
	13'h0cb5: q1 = 16'hd0bc; // 0x196a
	13'h0cb6: q1 = 16'h0000; // 0x196c
	13'h0cb7: q1 = 16'hcb8c; // 0x196e
	13'h0cb8: q1 = 16'h2040; // 0x1970
	13'h0cb9: q1 = 16'h1010; // 0x1972
	13'h0cba: q1 = 16'h4880; // 0x1974
	13'h0cbb: q1 = 16'h3740; // 0x1976
	13'h0cbc: q1 = 16'h0004; // 0x1978
	13'h0cbd: q1 = 16'h0c6b; // 0x197a
	13'h0cbe: q1 = 16'h0030; // 0x197c
	13'h0cbf: q1 = 16'h0004; // 0x197e
	13'h0cc0: q1 = 16'h670c; // 0x1980
	13'h0cc1: q1 = 16'h302b; // 0x1982
	13'h0cc2: q1 = 16'h0004; // 0x1984
	13'h0cc3: q1 = 16'h5240; // 0x1986
	13'h0cc4: q1 = 16'h3940; // 0x1988
	13'h0cc5: q1 = 16'h0014; // 0x198a
	13'h0cc6: q1 = 16'h600c; // 0x198c
	13'h0cc7: q1 = 16'h302c; // 0x198e
	13'h0cc8: q1 = 16'h0004; // 0x1990
	13'h0cc9: q1 = 16'hd07c; // 0x1992
	13'h0cca: q1 = 16'hffc0; // 0x1994
	13'h0ccb: q1 = 16'h3940; // 0x1996
	13'h0ccc: q1 = 16'h0014; // 0x1998
	13'h0ccd: q1 = 16'h302c; // 0x199a
	13'h0cce: q1 = 16'h0014; // 0x199c
	13'h0ccf: q1 = 16'h5240; // 0x199e
	13'h0cd0: q1 = 16'h3940; // 0x19a0
	13'h0cd1: q1 = 16'h001c; // 0x19a2
	13'h0cd2: q1 = 16'h397c; // 0x19a4
	13'h0cd3: q1 = 16'h000d; // 0x19a6
	13'h0cd4: q1 = 16'h000e; // 0x19a8
	13'h0cd5: q1 = 16'h377c; // 0x19aa
	13'h0cd6: q1 = 16'h001e; // 0x19ac
	13'h0cd7: q1 = 16'h0006; // 0x19ae
	13'h0cd8: q1 = 16'h397c; // 0x19b0
	13'h0cd9: q1 = 16'h001e; // 0x19b2
	13'h0cda: q1 = 16'h0016; // 0x19b4
	13'h0cdb: q1 = 16'h0c55; // 0x19b6
	13'h0cdc: q1 = 16'h0007; // 0x19b8
	13'h0cdd: q1 = 16'h6f0e; // 0x19ba
	13'h0cde: q1 = 16'h0c55; // 0x19bc
	13'h0cdf: q1 = 16'h000f; // 0x19be
	13'h0ce0: q1 = 16'h6c08; // 0x19c0
	13'h0ce1: q1 = 16'h397c; // 0x19c2
	13'h0ce2: q1 = 16'h001e; // 0x19c4
	13'h0ce3: q1 = 16'h001e; // 0x19c6
	13'h0ce4: q1 = 16'h6006; // 0x19c8
	13'h0ce5: q1 = 16'h397c; // 0x19ca
	13'h0ce6: q1 = 16'h000d; // 0x19cc
	13'h0ce7: q1 = 16'h001e; // 0x19ce
	13'h0ce8: q1 = 16'h206e; // 0x19d0
	13'h0ce9: q1 = 16'hfffc; // 0x19d2
	13'h0cea: q1 = 16'h317c; // 0x19d4
	13'h0ceb: q1 = 16'h0007; // 0x19d6
	13'h0cec: q1 = 16'h0006; // 0x19d8
	13'h0ced: q1 = 16'h206e; // 0x19da
	13'h0cee: q1 = 16'hfffc; // 0x19dc
	13'h0cef: q1 = 16'h3215; // 0x19de
	13'h0cf0: q1 = 16'h48c1; // 0x19e0
	13'h0cf1: q1 = 16'hd2bc; // 0x19e2
	13'h0cf2: q1 = 16'h0000; // 0x19e4
	13'h0cf3: q1 = 16'hcba4; // 0x19e6
	13'h0cf4: q1 = 16'h2241; // 0x19e8
	13'h0cf5: q1 = 16'h1211; // 0x19ea
	13'h0cf6: q1 = 16'h4881; // 0x19ec
	13'h0cf7: q1 = 16'h3141; // 0x19ee
	13'h0cf8: q1 = 16'h0004; // 0x19f0
	13'h0cf9: q1 = 16'h206e; // 0x19f2
	13'h0cfa: q1 = 16'hfffc; // 0x19f4
	13'h0cfb: q1 = 16'h3215; // 0x19f6
	13'h0cfc: q1 = 16'h48c1; // 0x19f8
	13'h0cfd: q1 = 16'hd2bc; // 0x19fa
	13'h0cfe: q1 = 16'h0000; // 0x19fc
	13'h0cff: q1 = 16'hcbbc; // 0x19fe
	13'h0d00: q1 = 16'h2241; // 0x1a00
	13'h0d01: q1 = 16'h1211; // 0x1a02
	13'h0d02: q1 = 16'h4881; // 0x1a04
	13'h0d03: q1 = 16'hef41; // 0x1a06
	13'h0d04: q1 = 16'hd254; // 0x1a08
	13'h0d05: q1 = 16'h3081; // 0x1a0a
	13'h0d06: q1 = 16'h206e; // 0x1a0c
	13'h0d07: q1 = 16'hfffc; // 0x1a0e
	13'h0d08: q1 = 16'h322c; // 0x1a10
	13'h0d09: q1 = 16'h0002; // 0x1a12
	13'h0d0a: q1 = 16'h3415; // 0x1a14
	13'h0d0b: q1 = 16'h48c2; // 0x1a16
	13'h0d0c: q1 = 16'hd4bc; // 0x1a18
	13'h0d0d: q1 = 16'h0000; // 0x1a1a
	13'h0d0e: q1 = 16'hcbd4; // 0x1a1c
	13'h0d0f: q1 = 16'h2442; // 0x1a1e
	13'h0d10: q1 = 16'h1412; // 0x1a20
	13'h0d11: q1 = 16'h4882; // 0x1a22
	13'h0d12: q1 = 16'hef42; // 0x1a24
	13'h0d13: q1 = 16'h9242; // 0x1a26
	13'h0d14: q1 = 16'h3141; // 0x1a28
	13'h0d15: q1 = 16'h0002; // 0x1a2a
	13'h0d16: q1 = 16'h0c55; // 0x1a2c
	13'h0d17: q1 = 16'h0014; // 0x1a2e
	13'h0d18: q1 = 16'h6c06; // 0x1a30
	13'h0d19: q1 = 16'h0c55; // 0x1a32
	13'h0d1a: q1 = 16'h0002; // 0x1a34
	13'h0d1b: q1 = 16'h6e2c; // 0x1a36
	13'h0d1c: q1 = 16'h7e02; // 0x1a38
	13'h0d1d: q1 = 16'h3007; // 0x1a3a
	13'h0d1e: q1 = 16'he740; // 0x1a3c
	13'h0d1f: q1 = 16'h48c0; // 0x1a3e
	13'h0d20: q1 = 16'h2840; // 0x1a40
	13'h0d21: q1 = 16'hd9fc; // 0x1a42
	13'h0d22: q1 = 16'h0001; // 0x1a44
	13'h0d23: q1 = 16'h8072; // 0x1a46
	13'h0d24: q1 = 16'hbe7c; // 0x1a48
	13'h0d25: q1 = 16'h0004; // 0x1a4a
	13'h0d26: q1 = 16'h6e16; // 0x1a4c
	13'h0d27: q1 = 16'h397c; // 0x1a4e
	13'h0d28: q1 = 16'h0030; // 0x1a50
	13'h0d29: q1 = 16'h0004; // 0x1a52
	13'h0d2a: q1 = 16'h426c; // 0x1a54
	13'h0d2b: q1 = 16'h0006; // 0x1a56
	13'h0d2c: q1 = 16'h4254; // 0x1a58
	13'h0d2d: q1 = 16'h426c; // 0x1a5a
	13'h0d2e: q1 = 16'h0002; // 0x1a5c
	13'h0d2f: q1 = 16'h5247; // 0x1a5e
	13'h0d30: q1 = 16'h508c; // 0x1a60
	13'h0d31: q1 = 16'h60e4; // 0x1a62
	13'h0d32: q1 = 16'h0c55; // 0x1a64
	13'h0d33: q1 = 16'h0013; // 0x1a66
	13'h0d34: q1 = 16'h6606; // 0x1a68
	13'h0d35: q1 = 16'h4eb9; // 0x1a6a
	13'h0d36: q1 = 16'h0000; // 0x1a6c
	13'h0d37: q1 = 16'h4162; // 0x1a6e
	13'h0d38: q1 = 16'h0c55; // 0x1a70
	13'h0d39: q1 = 16'h000f; // 0x1a72
	13'h0d3a: q1 = 16'h660c; // 0x1a74
	13'h0d3b: q1 = 16'h2ebc; // 0x1a76
	13'h0d3c: q1 = 16'h0000; // 0x1a78
	13'h0d3d: q1 = 16'hf6b0; // 0x1a7a
	13'h0d3e: q1 = 16'h4eb9; // 0x1a7c
	13'h0d3f: q1 = 16'h0000; // 0x1a7e
	13'h0d40: q1 = 16'h7dd8; // 0x1a80
	13'h0d41: q1 = 16'h0c55; // 0x1a82
	13'h0d42: q1 = 16'h000b; // 0x1a84
	13'h0d43: q1 = 16'h6d06; // 0x1a86
	13'h0d44: q1 = 16'h4eb9; // 0x1a88
	13'h0d45: q1 = 16'h0000; // 0x1a8a
	13'h0d46: q1 = 16'h4340; // 0x1a8c
	13'h0d47: q1 = 16'h5255; // 0x1a8e
	13'h0d48: q1 = 16'h4240; // 0x1a90
	13'h0d49: q1 = 16'h4a9f; // 0x1a92
	13'h0d4a: q1 = 16'h4cdf; // 0x1a94
	13'h0d4b: q1 = 16'h38c0; // 0x1a96
	13'h0d4c: q1 = 16'h4e5e; // 0x1a98
	13'h0d4d: q1 = 16'h4e75; // 0x1a9a
	13'h0d4e: q1 = 16'h4e56; // 0x1a9c
	13'h0d4f: q1 = 16'hfffc; // 0x1a9e
	13'h0d50: q1 = 16'h48e7; // 0x1aa0
	13'h0d51: q1 = 16'h0304; // 0x1aa2
	13'h0d52: q1 = 16'h2a7c; // 0x1aa4
	13'h0d53: q1 = 16'h0001; // 0x1aa6
	13'h0d54: q1 = 16'h7ec0; // 0x1aa8
	13'h0d55: q1 = 16'h4247; // 0x1aaa
	13'h0d56: q1 = 16'hbe7c; // 0x1aac
	13'h0d57: q1 = 16'h000a; // 0x1aae
	13'h0d58: q1 = 16'h6c1c; // 0x1ab0
	13'h0d59: q1 = 16'h4255; // 0x1ab2
	13'h0d5a: q1 = 16'h426d; // 0x1ab4
	13'h0d5b: q1 = 16'h0002; // 0x1ab6
	13'h0d5c: q1 = 16'h3007; // 0x1ab8
	13'h0d5d: q1 = 16'he540; // 0x1aba
	13'h0d5e: q1 = 16'h48c0; // 0x1abc
	13'h0d5f: q1 = 16'hd0bc; // 0x1abe
	13'h0d60: q1 = 16'h0001; // 0x1ac0
	13'h0d61: q1 = 16'h8902; // 0x1ac2
	13'h0d62: q1 = 16'h2040; // 0x1ac4
	13'h0d63: q1 = 16'h208d; // 0x1ac6
	13'h0d64: q1 = 16'h5c8d; // 0x1ac8
	13'h0d65: q1 = 16'h5247; // 0x1aca
	13'h0d66: q1 = 16'h60de; // 0x1acc
	13'h0d67: q1 = 16'h2079; // 0x1ace
	13'h0d68: q1 = 16'h0001; // 0x1ad0
	13'h0d69: q1 = 16'h7fb8; // 0x1ad2
	13'h0d6a: q1 = 16'h3010; // 0x1ad4
	13'h0d6b: q1 = 16'h5440; // 0x1ad6
	13'h0d6c: q1 = 16'h33c0; // 0x1ad8
	13'h0d6d: q1 = 16'h0001; // 0x1ada
	13'h0d6e: q1 = 16'h7fd2; // 0x1adc
	13'h0d6f: q1 = 16'h0c79; // 0x1ade
	13'h0d70: q1 = 16'h000a; // 0x1ae0
	13'h0d71: q1 = 16'h0001; // 0x1ae2
	13'h0d72: q1 = 16'h7fd2; // 0x1ae4
	13'h0d73: q1 = 16'h6f08; // 0x1ae6
	13'h0d74: q1 = 16'h33fc; // 0x1ae8
	13'h0d75: q1 = 16'h000a; // 0x1aea
	13'h0d76: q1 = 16'h0001; // 0x1aec
	13'h0d77: q1 = 16'h7fd2; // 0x1aee
	13'h0d78: q1 = 16'h2a7c; // 0x1af0
	13'h0d79: q1 = 16'h0001; // 0x1af2
	13'h0d7a: q1 = 16'h7ec0; // 0x1af4
	13'h0d7b: q1 = 16'h4247; // 0x1af6
	13'h0d7c: q1 = 16'hbe79; // 0x1af8
	13'h0d7d: q1 = 16'h0001; // 0x1afa
	13'h0d7e: q1 = 16'h7fd2; // 0x1afc
	13'h0d7f: q1 = 16'h6c00; // 0x1afe
	13'h0d80: q1 = 16'h00d6; // 0x1b00
	13'h0d81: q1 = 16'h3ebc; // 0x1b02
	13'h0d82: q1 = 16'h7700; // 0x1b04
	13'h0d83: q1 = 16'h3f3c; // 0x1b06
	13'h0d84: q1 = 16'h0580; // 0x1b08
	13'h0d85: q1 = 16'h4eb9; // 0x1b0a
	13'h0d86: q1 = 16'h0000; // 0x1b0c
	13'h0d87: q1 = 16'h8e6c; // 0x1b0e
	13'h0d88: q1 = 16'h4a5f; // 0x1b10
	13'h0d89: q1 = 16'h3d40; // 0x1b12
	13'h0d8a: q1 = 16'hfffe; // 0x1b14
	13'h0d8b: q1 = 16'h3ebc; // 0x1b16
	13'h0d8c: q1 = 16'h7380; // 0x1b18
	13'h0d8d: q1 = 16'h3f3c; // 0x1b1a
	13'h0d8e: q1 = 16'h1800; // 0x1b1c
	13'h0d8f: q1 = 16'h4eb9; // 0x1b1e
	13'h0d90: q1 = 16'h0000; // 0x1b20
	13'h0d91: q1 = 16'h8e6c; // 0x1b22
	13'h0d92: q1 = 16'h4a5f; // 0x1b24
	13'h0d93: q1 = 16'h3d40; // 0x1b26
	13'h0d94: q1 = 16'hfffc; // 0x1b28
	13'h0d95: q1 = 16'h200e; // 0x1b2a
	13'h0d96: q1 = 16'hd0bc; // 0x1b2c
	13'h0d97: q1 = 16'hffff; // 0x1b2e
	13'h0d98: q1 = 16'hfffc; // 0x1b30
	13'h0d99: q1 = 16'h2e80; // 0x1b32
	13'h0d9a: q1 = 16'h200e; // 0x1b34
	13'h0d9b: q1 = 16'hd0bc; // 0x1b36
	13'h0d9c: q1 = 16'hffff; // 0x1b38
	13'h0d9d: q1 = 16'hfffe; // 0x1b3a
	13'h0d9e: q1 = 16'h2f00; // 0x1b3c
	13'h0d9f: q1 = 16'h4eb9; // 0x1b3e
	13'h0da0: q1 = 16'h0000; // 0x1b40
	13'h0da1: q1 = 16'hbee0; // 0x1b42
	13'h0da2: q1 = 16'h4a9f; // 0x1b44
	13'h0da3: q1 = 16'h3eae; // 0x1b46
	13'h0da4: q1 = 16'hfffc; // 0x1b48
	13'h0da5: q1 = 16'h3f2e; // 0x1b4a
	13'h0da6: q1 = 16'hfffe; // 0x1b4c
	13'h0da7: q1 = 16'h4eb9; // 0x1b4e
	13'h0da8: q1 = 16'h0000; // 0x1b50
	13'h0da9: q1 = 16'h4d7e; // 0x1b52
	13'h0daa: q1 = 16'h4a5f; // 0x1b54
	13'h0dab: q1 = 16'h4a40; // 0x1b56
	13'h0dac: q1 = 16'h66a8; // 0x1b58
	13'h0dad: q1 = 16'h3ebc; // 0x1b5a
	13'h0dae: q1 = 16'h0001; // 0x1b5c
	13'h0daf: q1 = 16'h200e; // 0x1b5e
	13'h0db0: q1 = 16'hd0bc; // 0x1b60
	13'h0db1: q1 = 16'hffff; // 0x1b62
	13'h0db2: q1 = 16'hfffc; // 0x1b64
	13'h0db3: q1 = 16'h2f00; // 0x1b66
	13'h0db4: q1 = 16'h200e; // 0x1b68
	13'h0db5: q1 = 16'hd0bc; // 0x1b6a
	13'h0db6: q1 = 16'hffff; // 0x1b6c
	13'h0db7: q1 = 16'hfffe; // 0x1b6e
	13'h0db8: q1 = 16'h2f00; // 0x1b70
	13'h0db9: q1 = 16'h4eb9; // 0x1b72
	13'h0dba: q1 = 16'h0000; // 0x1b74
	13'h0dbb: q1 = 16'h5d44; // 0x1b76
	13'h0dbc: q1 = 16'hbf8f; // 0x1b78
	13'h0dbd: q1 = 16'h4a40; // 0x1b7a
	13'h0dbe: q1 = 16'h6684; // 0x1b7c
	13'h0dbf: q1 = 16'h3ebc; // 0x1b7e
	13'h0dc0: q1 = 16'h0001; // 0x1b80
	13'h0dc1: q1 = 16'h3f2e; // 0x1b82
	13'h0dc2: q1 = 16'hfffc; // 0x1b84
	13'h0dc3: q1 = 16'h3f2e; // 0x1b86
	13'h0dc4: q1 = 16'hfffe; // 0x1b88
	13'h0dc5: q1 = 16'h4eb9; // 0x1b8a
	13'h0dc6: q1 = 16'h0000; // 0x1b8c
	13'h0dc7: q1 = 16'h8744; // 0x1b8e
	13'h0dc8: q1 = 16'h4a9f; // 0x1b90
	13'h0dc9: q1 = 16'h4a40; // 0x1b92
	13'h0dca: q1 = 16'h6600; // 0x1b94
	13'h0dcb: q1 = 16'hff6c; // 0x1b96
	13'h0dcc: q1 = 16'h3ebc; // 0x1b98
	13'h0dcd: q1 = 16'h0001; // 0x1b9a
	13'h0dce: q1 = 16'h3f2e; // 0x1b9c
	13'h0dcf: q1 = 16'hfffc; // 0x1b9e
	13'h0dd0: q1 = 16'h3f2e; // 0x1ba0
	13'h0dd1: q1 = 16'hfffe; // 0x1ba2
	13'h0dd2: q1 = 16'h4eb9; // 0x1ba4
	13'h0dd3: q1 = 16'h0000; // 0x1ba6
	13'h0dd4: q1 = 16'h42d4; // 0x1ba8
	13'h0dd5: q1 = 16'h4a9f; // 0x1baa
	13'h0dd6: q1 = 16'h4a40; // 0x1bac
	13'h0dd7: q1 = 16'h6600; // 0x1bae
	13'h0dd8: q1 = 16'hff52; // 0x1bb0
	13'h0dd9: q1 = 16'h6004; // 0x1bb2
	13'h0dda: q1 = 16'h6000; // 0x1bb4
	13'h0ddb: q1 = 16'hff4c; // 0x1bb6
	13'h0ddc: q1 = 16'h3aae; // 0x1bb8
	13'h0ddd: q1 = 16'hfffe; // 0x1bba
	13'h0dde: q1 = 16'h3b6e; // 0x1bbc
	13'h0ddf: q1 = 16'hfffc; // 0x1bbe
	13'h0de0: q1 = 16'h0002; // 0x1bc0
	13'h0de1: q1 = 16'h4257; // 0x1bc2
	13'h0de2: q1 = 16'h2f0d; // 0x1bc4
	13'h0de3: q1 = 16'h4eb9; // 0x1bc6
	13'h0de4: q1 = 16'h0000; // 0x1bc8
	13'h0de5: q1 = 16'h5f04; // 0x1bca
	13'h0de6: q1 = 16'h4a9f; // 0x1bcc
	13'h0de7: q1 = 16'h5c8d; // 0x1bce
	13'h0de8: q1 = 16'h5247; // 0x1bd0
	13'h0de9: q1 = 16'h6000; // 0x1bd2
	13'h0dea: q1 = 16'hff24; // 0x1bd4
	13'h0deb: q1 = 16'h4a9f; // 0x1bd6
	13'h0dec: q1 = 16'h4cdf; // 0x1bd8
	13'h0ded: q1 = 16'h2080; // 0x1bda
	13'h0dee: q1 = 16'h4e5e; // 0x1bdc
	13'h0def: q1 = 16'h4e75; // 0x1bde
	13'h0df0: q1 = 16'h4e56; // 0x1be0
	13'h0df1: q1 = 16'hfff4; // 0x1be2
	13'h0df2: q1 = 16'h48e7; // 0x1be4
	13'h0df3: q1 = 16'h0704; // 0x1be6
	13'h0df4: q1 = 16'h4a6e; // 0x1be8
	13'h0df5: q1 = 16'h0008; // 0x1bea
	13'h0df6: q1 = 16'h6646; // 0x1bec
	13'h0df7: q1 = 16'h33fc; // 0x1bee
	13'h0df8: q1 = 16'h0004; // 0x1bf0
	13'h0df9: q1 = 16'h0001; // 0x1bf2
	13'h0dfa: q1 = 16'h7fd2; // 0x1bf4
	13'h0dfb: q1 = 16'h2a7c; // 0x1bf6
	13'h0dfc: q1 = 16'h0001; // 0x1bf8
	13'h0dfd: q1 = 16'h7ec0; // 0x1bfa
	13'h0dfe: q1 = 16'h4247; // 0x1bfc
	13'h0dff: q1 = 16'hbe79; // 0x1bfe
	13'h0e00: q1 = 16'h0001; // 0x1c00
	13'h0e01: q1 = 16'h7fd2; // 0x1c02
	13'h0e02: q1 = 16'h6c2a; // 0x1c04
	13'h0e03: q1 = 16'h3abc; // 0x1c06
	13'h0e04: q1 = 16'h0800; // 0x1c08
	13'h0e05: q1 = 16'h7014; // 0x1c0a
	13'h0e06: q1 = 16'h3207; // 0x1c0c
	13'h0e07: q1 = 16'hc3fc; // 0x1c0e
	13'h0e08: q1 = 16'h0003; // 0x1c10
	13'h0e09: q1 = 16'h9041; // 0x1c12
	13'h0e0a: q1 = 16'h4281; // 0x1c14
	13'h0e0b: q1 = 16'h720a; // 0x1c16
	13'h0e0c: q1 = 16'he360; // 0x1c18
	13'h0e0d: q1 = 16'h3b40; // 0x1c1a
	13'h0e0e: q1 = 16'h0002; // 0x1c1c
	13'h0e0f: q1 = 16'h4257; // 0x1c1e
	13'h0e10: q1 = 16'h2f0d; // 0x1c20
	13'h0e11: q1 = 16'h4eb9; // 0x1c22
	13'h0e12: q1 = 16'h0000; // 0x1c24
	13'h0e13: q1 = 16'h5f04; // 0x1c26
	13'h0e14: q1 = 16'h4a9f; // 0x1c28
	13'h0e15: q1 = 16'h5c8d; // 0x1c2a
	13'h0e16: q1 = 16'h5247; // 0x1c2c
	13'h0e17: q1 = 16'h60ce; // 0x1c2e
	13'h0e18: q1 = 16'h6000; // 0x1c30
	13'h0e19: q1 = 16'h0108; // 0x1c32
	13'h0e1a: q1 = 16'h0c6e; // 0x1c34
	13'h0e1b: q1 = 16'h0002; // 0x1c36
	13'h0e1c: q1 = 16'h0008; // 0x1c38
	13'h0e1d: q1 = 16'h660a; // 0x1c3a
	13'h0e1e: q1 = 16'h4279; // 0x1c3c
	13'h0e1f: q1 = 16'h0001; // 0x1c3e
	13'h0e20: q1 = 16'h7fd2; // 0x1c40
	13'h0e21: q1 = 16'h6000; // 0x1c42
	13'h0e22: q1 = 16'h00f6; // 0x1c44
	13'h0e23: q1 = 16'h0c6e; // 0x1c46
	13'h0e24: q1 = 16'h0003; // 0x1c48
	13'h0e25: q1 = 16'h0008; // 0x1c4a
	13'h0e26: q1 = 16'h6660; // 0x1c4c
	13'h0e27: q1 = 16'h33fc; // 0x1c4e
	13'h0e28: q1 = 16'h0005; // 0x1c50
	13'h0e29: q1 = 16'h0001; // 0x1c52
	13'h0e2a: q1 = 16'h7fd2; // 0x1c54
	13'h0e2b: q1 = 16'h2a7c; // 0x1c56
	13'h0e2c: q1 = 16'h0001; // 0x1c58
	13'h0e2d: q1 = 16'h7ec0; // 0x1c5a
	13'h0e2e: q1 = 16'h4247; // 0x1c5c
	13'h0e2f: q1 = 16'hbe79; // 0x1c5e
	13'h0e30: q1 = 16'h0001; // 0x1c60
	13'h0e31: q1 = 16'h7fd2; // 0x1c62
	13'h0e32: q1 = 16'h6c44; // 0x1c64
	13'h0e33: q1 = 16'h3007; // 0x1c66
	13'h0e34: q1 = 16'he340; // 0x1c68
	13'h0e35: q1 = 16'h48c0; // 0x1c6a
	13'h0e36: q1 = 16'hd0bc; // 0x1c6c
	13'h0e37: q1 = 16'h0000; // 0x1c6e
	13'h0e38: q1 = 16'hcc1c; // 0x1c70
	13'h0e39: q1 = 16'h2040; // 0x1c72
	13'h0e3a: q1 = 16'h3010; // 0x1c74
	13'h0e3b: q1 = 16'h4281; // 0x1c76
	13'h0e3c: q1 = 16'h720a; // 0x1c78
	13'h0e3d: q1 = 16'he360; // 0x1c7a
	13'h0e3e: q1 = 16'h3a80; // 0x1c7c
	13'h0e3f: q1 = 16'h3007; // 0x1c7e
	13'h0e40: q1 = 16'he340; // 0x1c80
	13'h0e41: q1 = 16'h48c0; // 0x1c82
	13'h0e42: q1 = 16'hd0bc; // 0x1c84
	13'h0e43: q1 = 16'h0000; // 0x1c86
	13'h0e44: q1 = 16'hcc26; // 0x1c88
	13'h0e45: q1 = 16'h2040; // 0x1c8a
	13'h0e46: q1 = 16'h3010; // 0x1c8c
	13'h0e47: q1 = 16'h4281; // 0x1c8e
	13'h0e48: q1 = 16'h720a; // 0x1c90
	13'h0e49: q1 = 16'he360; // 0x1c92
	13'h0e4a: q1 = 16'h3b40; // 0x1c94
	13'h0e4b: q1 = 16'h0002; // 0x1c96
	13'h0e4c: q1 = 16'h4257; // 0x1c98
	13'h0e4d: q1 = 16'h2f0d; // 0x1c9a
	13'h0e4e: q1 = 16'h4eb9; // 0x1c9c
	13'h0e4f: q1 = 16'h0000; // 0x1c9e
	13'h0e50: q1 = 16'h5f04; // 0x1ca0
	13'h0e51: q1 = 16'h4a9f; // 0x1ca2
	13'h0e52: q1 = 16'h5c8d; // 0x1ca4
	13'h0e53: q1 = 16'h5247; // 0x1ca6
	13'h0e54: q1 = 16'h60b4; // 0x1ca8
	13'h0e55: q1 = 16'h6000; // 0x1caa
	13'h0e56: q1 = 16'h008e; // 0x1cac
	13'h0e57: q1 = 16'h0c6e; // 0x1cae
	13'h0e58: q1 = 16'h0006; // 0x1cb0
	13'h0e59: q1 = 16'h0008; // 0x1cb2
	13'h0e5a: q1 = 16'h670a; // 0x1cb4
	13'h0e5b: q1 = 16'h0c6e; // 0x1cb6
	13'h0e5c: q1 = 16'h0007; // 0x1cb8
	13'h0e5d: q1 = 16'h0008; // 0x1cba
	13'h0e5e: q1 = 16'h6600; // 0x1cbc
	13'h0e5f: q1 = 16'h007c; // 0x1cbe
	13'h0e60: q1 = 16'h0c6e; // 0x1cc0
	13'h0e61: q1 = 16'h0006; // 0x1cc2
	13'h0e62: q1 = 16'h0008; // 0x1cc4
	13'h0e63: q1 = 16'h6604; // 0x1cc6
	13'h0e64: q1 = 16'h7c3e; // 0x1cc8
	13'h0e65: q1 = 16'h6002; // 0x1cca
	13'h0e66: q1 = 16'h4246; // 0x1ccc
	13'h0e67: q1 = 16'h3ebc; // 0x1cce
	13'h0e68: q1 = 16'h002f; // 0x1cd0
	13'h0e69: q1 = 16'h200e; // 0x1cd2
	13'h0e6a: q1 = 16'hd0bc; // 0x1cd4
	13'h0e6b: q1 = 16'hffff; // 0x1cd6
	13'h0e6c: q1 = 16'hfff4; // 0x1cd8
	13'h0e6d: q1 = 16'h2f00; // 0x1cda
	13'h0e6e: q1 = 16'h4eb9; // 0x1cdc
	13'h0e6f: q1 = 16'h0000; // 0x1cde
	13'h0e70: q1 = 16'h78f6; // 0x1ce0
	13'h0e71: q1 = 16'h4a9f; // 0x1ce2
	13'h0e72: q1 = 16'h3e86; // 0x1ce4
	13'h0e73: q1 = 16'h4267; // 0x1ce6
	13'h0e74: q1 = 16'h3f3c; // 0x1ce8
	13'h0e75: q1 = 16'h0007; // 0x1cea
	13'h0e76: q1 = 16'h3f3c; // 0x1cec
	13'h0e77: q1 = 16'h000f; // 0x1cee
	13'h0e78: q1 = 16'h200e; // 0x1cf0
	13'h0e79: q1 = 16'hd0bc; // 0x1cf2
	13'h0e7a: q1 = 16'hffff; // 0x1cf4
	13'h0e7b: q1 = 16'hfff4; // 0x1cf6
	13'h0e7c: q1 = 16'h2f00; // 0x1cf8
	13'h0e7d: q1 = 16'h4eb9; // 0x1cfa
	13'h0e7e: q1 = 16'h0000; // 0x1cfc
	13'h0e7f: q1 = 16'h026c; // 0x1cfe
	13'h0e80: q1 = 16'hdefc; // 0x1d00
	13'h0e81: q1 = 16'h000a; // 0x1d02
	13'h0e82: q1 = 16'h3ebc; // 0x1d04
	13'h0e83: q1 = 16'h0030; // 0x1d06
	13'h0e84: q1 = 16'h200e; // 0x1d08
	13'h0e85: q1 = 16'hd0bc; // 0x1d0a
	13'h0e86: q1 = 16'hffff; // 0x1d0c
	13'h0e87: q1 = 16'hfff4; // 0x1d0e
	13'h0e88: q1 = 16'h2f00; // 0x1d10
	13'h0e89: q1 = 16'h4eb9; // 0x1d12
	13'h0e8a: q1 = 16'h0000; // 0x1d14
	13'h0e8b: q1 = 16'h78f6; // 0x1d16
	13'h0e8c: q1 = 16'h4a9f; // 0x1d18
	13'h0e8d: q1 = 16'h3e86; // 0x1d1a
	13'h0e8e: q1 = 16'h4267; // 0x1d1c
	13'h0e8f: q1 = 16'h3f3c; // 0x1d1e
	13'h0e90: q1 = 16'h0009; // 0x1d20
	13'h0e91: q1 = 16'h3f3c; // 0x1d22
	13'h0e92: q1 = 16'h000c; // 0x1d24
	13'h0e93: q1 = 16'h200e; // 0x1d26
	13'h0e94: q1 = 16'hd0bc; // 0x1d28
	13'h0e95: q1 = 16'hffff; // 0x1d2a
	13'h0e96: q1 = 16'hfff4; // 0x1d2c
	13'h0e97: q1 = 16'h2f00; // 0x1d2e
	13'h0e98: q1 = 16'h4eb9; // 0x1d30
	13'h0e99: q1 = 16'h0000; // 0x1d32
	13'h0e9a: q1 = 16'h026c; // 0x1d34
	13'h0e9b: q1 = 16'hdefc; // 0x1d36
	13'h0e9c: q1 = 16'h000a; // 0x1d38
	13'h0e9d: q1 = 16'h4a9f; // 0x1d3a
	13'h0e9e: q1 = 16'h4cdf; // 0x1d3c
	13'h0e9f: q1 = 16'h20c0; // 0x1d3e
	13'h0ea0: q1 = 16'h4e5e; // 0x1d40
	13'h0ea1: q1 = 16'h4e75; // 0x1d42
	13'h0ea2: q1 = 16'h4e56; // 0x1d44
	13'h0ea3: q1 = 16'hfffc; // 0x1d46
	13'h0ea4: q1 = 16'h48e7; // 0x1d48
	13'h0ea5: q1 = 16'h0f1c; // 0x1d4a
	13'h0ea6: q1 = 16'h2a6e; // 0x1d4c
	13'h0ea7: q1 = 16'h0008; // 0x1d4e
	13'h0ea8: q1 = 16'h286e; // 0x1d50
	13'h0ea9: q1 = 16'h000c; // 0x1d52
	13'h0eaa: q1 = 16'h3e2e; // 0x1d54
	13'h0eab: q1 = 16'h0010; // 0x1d56
	13'h0eac: q1 = 16'hbe7c; // 0x1d58
	13'h0ead: q1 = 16'h0001; // 0x1d5a
	13'h0eae: q1 = 16'h6670; // 0x1d5c
	13'h0eaf: q1 = 16'h3d7c; // 0x1d5e
	13'h0eb0: q1 = 16'h1000; // 0x1d60
	13'h0eb1: q1 = 16'hfffe; // 0x1d62
	13'h0eb2: q1 = 16'h3d7c; // 0x1d64
	13'h0eb3: q1 = 16'h1000; // 0x1d66
	13'h0eb4: q1 = 16'hfffc; // 0x1d68
	13'h0eb5: q1 = 16'h0c79; // 0x1d6a
	13'h0eb6: q1 = 16'h0006; // 0x1d6c
	13'h0eb7: q1 = 16'h0001; // 0x1d6e
	13'h0eb8: q1 = 16'h7fd2; // 0x1d70
	13'h0eb9: q1 = 16'h6d06; // 0x1d72
	13'h0eba: q1 = 16'h3d7c; // 0x1d74
	13'h0ebb: q1 = 16'h0c00; // 0x1d76
	13'h0ebc: q1 = 16'hfffe; // 0x1d78
	13'h0ebd: q1 = 16'h0c79; // 0x1d7a
	13'h0ebe: q1 = 16'h0008; // 0x1d7c
	13'h0ebf: q1 = 16'h0001; // 0x1d7e
	13'h0ec0: q1 = 16'h7fd2; // 0x1d80
	13'h0ec1: q1 = 16'h6d06; // 0x1d82
	13'h0ec2: q1 = 16'h3d7c; // 0x1d84
	13'h0ec3: q1 = 16'h0800; // 0x1d86
	13'h0ec4: q1 = 16'hfffc; // 0x1d88
	13'h0ec5: q1 = 16'h267c; // 0x1d8a
	13'h0ec6: q1 = 16'h0001; // 0x1d8c
	13'h0ec7: q1 = 16'h7ec0; // 0x1d8e
	13'h0ec8: q1 = 16'h4246; // 0x1d90
	13'h0ec9: q1 = 16'hbc79; // 0x1d92
	13'h0eca: q1 = 16'h0001; // 0x1d94
	13'h0ecb: q1 = 16'h7fd2; // 0x1d96
	13'h0ecc: q1 = 16'h6c32; // 0x1d98
	13'h0ecd: q1 = 16'h3e95; // 0x1d9a
	13'h0ece: q1 = 16'h3013; // 0x1d9c
	13'h0ecf: q1 = 16'h9157; // 0x1d9e
	13'h0ed0: q1 = 16'h4eb9; // 0x1da0
	13'h0ed1: q1 = 16'h0000; // 0x1da2
	13'h0ed2: q1 = 16'h09a2; // 0x1da4
	13'h0ed3: q1 = 16'hb06e; // 0x1da6
	13'h0ed4: q1 = 16'hfffe; // 0x1da8
	13'h0ed5: q1 = 16'h6c1a; // 0x1daa
	13'h0ed6: q1 = 16'h3e94; // 0x1dac
	13'h0ed7: q1 = 16'h302b; // 0x1dae
	13'h0ed8: q1 = 16'h0002; // 0x1db0
	13'h0ed9: q1 = 16'h9157; // 0x1db2
	13'h0eda: q1 = 16'h4eb9; // 0x1db4
	13'h0edb: q1 = 16'h0000; // 0x1db6
	13'h0edc: q1 = 16'h09a2; // 0x1db8
	13'h0edd: q1 = 16'hb06e; // 0x1dba
	13'h0ede: q1 = 16'hfffc; // 0x1dbc
	13'h0edf: q1 = 16'h6c06; // 0x1dbe
	13'h0ee0: q1 = 16'h7001; // 0x1dc0
	13'h0ee1: q1 = 16'h6000; // 0x1dc2
	13'h0ee2: q1 = 16'h006c; // 0x1dc4
	13'h0ee3: q1 = 16'h5c8b; // 0x1dc6
	13'h0ee4: q1 = 16'h5246; // 0x1dc8
	13'h0ee5: q1 = 16'h60c6; // 0x1dca
	13'h0ee6: q1 = 16'h6060; // 0x1dcc
	13'h0ee7: q1 = 16'h267c; // 0x1dce
	13'h0ee8: q1 = 16'h0001; // 0x1dd0
	13'h0ee9: q1 = 16'h7ec0; // 0x1dd2
	13'h0eea: q1 = 16'h4246; // 0x1dd4
	13'h0eeb: q1 = 16'hbc79; // 0x1dd6
	13'h0eec: q1 = 16'h0001; // 0x1dd8
	13'h0eed: q1 = 16'h7fd2; // 0x1dda
	13'h0eee: q1 = 16'h6c50; // 0x1ddc
	13'h0eef: q1 = 16'h0c6b; // 0x1dde
	13'h0ef0: q1 = 16'h0001; // 0x1de0
	13'h0ef1: q1 = 16'h0004; // 0x1de2
	13'h0ef2: q1 = 16'h6642; // 0x1de4
	13'h0ef3: q1 = 16'h3a15; // 0x1de6
	13'h0ef4: q1 = 16'h9a53; // 0x1de8
	13'h0ef5: q1 = 16'h4a45; // 0x1dea
	13'h0ef6: q1 = 16'h6c06; // 0x1dec
	13'h0ef7: q1 = 16'h3005; // 0x1dee
	13'h0ef8: q1 = 16'h4440; // 0x1df0
	13'h0ef9: q1 = 16'h3a00; // 0x1df2
	13'h0efa: q1 = 16'hba7c; // 0x1df4
	13'h0efb: q1 = 16'h0500; // 0x1df6
	13'h0efc: q1 = 16'h6c2e; // 0x1df8
	13'h0efd: q1 = 16'h3014; // 0x1dfa
	13'h0efe: q1 = 16'h322b; // 0x1dfc
	13'h0eff: q1 = 16'h0002; // 0x1dfe
	13'h0f00: q1 = 16'hd27c; // 0x1e00
	13'h0f01: q1 = 16'h0100; // 0x1e02
	13'h0f02: q1 = 16'h9041; // 0x1e04
	13'h0f03: q1 = 16'h3a00; // 0x1e06
	13'h0f04: q1 = 16'h4a45; // 0x1e08
	13'h0f05: q1 = 16'h6c06; // 0x1e0a
	13'h0f06: q1 = 16'h3005; // 0x1e0c
	13'h0f07: q1 = 16'h4440; // 0x1e0e
	13'h0f08: q1 = 16'h3a00; // 0x1e10
	13'h0f09: q1 = 16'hba7c; // 0x1e12
	13'h0f0a: q1 = 16'h0200; // 0x1e14
	13'h0f0b: q1 = 16'h6c10; // 0x1e16
	13'h0f0c: q1 = 16'h3a93; // 0x1e18
	13'h0f0d: q1 = 16'h302b; // 0x1e1a
	13'h0f0e: q1 = 16'h0002; // 0x1e1c
	13'h0f0f: q1 = 16'hd07c; // 0x1e1e
	13'h0f10: q1 = 16'h0100; // 0x1e20
	13'h0f11: q1 = 16'h3880; // 0x1e22
	13'h0f12: q1 = 16'h7001; // 0x1e24
	13'h0f13: q1 = 16'h6008; // 0x1e26
	13'h0f14: q1 = 16'h5c8b; // 0x1e28
	13'h0f15: q1 = 16'h5246; // 0x1e2a
	13'h0f16: q1 = 16'h60a8; // 0x1e2c
	13'h0f17: q1 = 16'h4240; // 0x1e2e
	13'h0f18: q1 = 16'h4a9f; // 0x1e30
	13'h0f19: q1 = 16'h4cdf; // 0x1e32
	13'h0f1a: q1 = 16'h38e0; // 0x1e34
	13'h0f1b: q1 = 16'h4e5e; // 0x1e36
	13'h0f1c: q1 = 16'h4e75; // 0x1e38
	13'h0f1d: q1 = 16'h4e56; // 0x1e3a
	13'h0f1e: q1 = 16'h0000; // 0x1e3c
	13'h0f1f: q1 = 16'h48e7; // 0x1e3e
	13'h0f20: q1 = 16'h0304; // 0x1e40
	13'h0f21: q1 = 16'h4a6e; // 0x1e42
	13'h0f22: q1 = 16'h0010; // 0x1e44
	13'h0f23: q1 = 16'h6630; // 0x1e46
	13'h0f24: q1 = 16'h3eb9; // 0x1e48
	13'h0f25: q1 = 16'h0001; // 0x1e4a
	13'h0f26: q1 = 16'h7fd2; // 0x1e4c
	13'h0f27: q1 = 16'h5357; // 0x1e4e
	13'h0f28: q1 = 16'h4267; // 0x1e50
	13'h0f29: q1 = 16'h4eb9; // 0x1e52
	13'h0f2a: q1 = 16'h0000; // 0x1e54
	13'h0f2b: q1 = 16'h8e6c; // 0x1e56
	13'h0f2c: q1 = 16'h4a5f; // 0x1e58
	13'h0f2d: q1 = 16'h3e00; // 0x1e5a
	13'h0f2e: q1 = 16'h3007; // 0x1e5c
	13'h0f2f: q1 = 16'he540; // 0x1e5e
	13'h0f30: q1 = 16'h48c0; // 0x1e60
	13'h0f31: q1 = 16'hd0bc; // 0x1e62
	13'h0f32: q1 = 16'h0001; // 0x1e64
	13'h0f33: q1 = 16'h8902; // 0x1e66
	13'h0f34: q1 = 16'h2040; // 0x1e68
	13'h0f35: q1 = 16'h2a50; // 0x1e6a
	13'h0f36: q1 = 16'h0c6d; // 0x1e6c
	13'h0f37: q1 = 16'h0002; // 0x1e6e
	13'h0f38: q1 = 16'h0004; // 0x1e70
	13'h0f39: q1 = 16'h6602; // 0x1e72
	13'h0f3a: q1 = 16'h60d2; // 0x1e74
	13'h0f3b: q1 = 16'h6014; // 0x1e76
	13'h0f3c: q1 = 16'h302e; // 0x1e78
	13'h0f3d: q1 = 16'h0010; // 0x1e7a
	13'h0f3e: q1 = 16'h5340; // 0x1e7c
	13'h0f3f: q1 = 16'he540; // 0x1e7e
	13'h0f40: q1 = 16'h48c0; // 0x1e80
	13'h0f41: q1 = 16'hd0bc; // 0x1e82
	13'h0f42: q1 = 16'h0001; // 0x1e84
	13'h0f43: q1 = 16'h8902; // 0x1e86
	13'h0f44: q1 = 16'h2040; // 0x1e88
	13'h0f45: q1 = 16'h2a50; // 0x1e8a
	13'h0f46: q1 = 16'h206e; // 0x1e8c
	13'h0f47: q1 = 16'h0008; // 0x1e8e
	13'h0f48: q1 = 16'h3095; // 0x1e90
	13'h0f49: q1 = 16'h206e; // 0x1e92
	13'h0f4a: q1 = 16'h000c; // 0x1e94
	13'h0f4b: q1 = 16'h322d; // 0x1e96
	13'h0f4c: q1 = 16'h0002; // 0x1e98
	13'h0f4d: q1 = 16'hd27c; // 0x1e9a
	13'h0f4e: q1 = 16'h0100; // 0x1e9c
	13'h0f4f: q1 = 16'h3081; // 0x1e9e
	13'h0f50: q1 = 16'h3b7c; // 0x1ea0
	13'h0f51: q1 = 16'h0002; // 0x1ea2
	13'h0f52: q1 = 16'h0004; // 0x1ea4
	13'h0f53: q1 = 16'h4a9f; // 0x1ea6
	13'h0f54: q1 = 16'h4cdf; // 0x1ea8
	13'h0f55: q1 = 16'h2080; // 0x1eaa
	13'h0f56: q1 = 16'h4e5e; // 0x1eac
	13'h0f57: q1 = 16'h4e75; // 0x1eae
	13'h0f58: q1 = 16'h4e56; // 0x1eb0
	13'h0f59: q1 = 16'h0000; // 0x1eb2
	13'h0f5a: q1 = 16'h48e7; // 0x1eb4
	13'h0f5b: q1 = 16'h0304; // 0x1eb6
	13'h0f5c: q1 = 16'h4247; // 0x1eb8
	13'h0f5d: q1 = 16'h2a7c; // 0x1eba
	13'h0f5e: q1 = 16'h0001; // 0x1ebc
	13'h0f5f: q1 = 16'h7ec0; // 0x1ebe
	13'h0f60: q1 = 16'hbe79; // 0x1ec0
	13'h0f61: q1 = 16'h0001; // 0x1ec2
	13'h0f62: q1 = 16'h7fd2; // 0x1ec4
	13'h0f63: q1 = 16'h6c1c; // 0x1ec6
	13'h0f64: q1 = 16'h3015; // 0x1ec8
	13'h0f65: q1 = 16'hb06e; // 0x1eca
	13'h0f66: q1 = 16'h0008; // 0x1ecc
	13'h0f67: q1 = 16'h660e; // 0x1ece
	13'h0f68: q1 = 16'h302e; // 0x1ed0
	13'h0f69: q1 = 16'h000a; // 0x1ed2
	13'h0f6a: q1 = 16'hd07c; // 0x1ed4
	13'h0f6b: q1 = 16'hff00; // 0x1ed6
	13'h0f6c: q1 = 16'hb06d; // 0x1ed8
	13'h0f6d: q1 = 16'h0002; // 0x1eda
	13'h0f6e: q1 = 16'h6706; // 0x1edc
	13'h0f6f: q1 = 16'h5c8d; // 0x1ede
	13'h0f70: q1 = 16'h5247; // 0x1ee0
	13'h0f71: q1 = 16'h60dc; // 0x1ee2
	13'h0f72: q1 = 16'hbe79; // 0x1ee4
	13'h0f73: q1 = 16'h0001; // 0x1ee6
	13'h0f74: q1 = 16'h7fd2; // 0x1ee8
	13'h0f75: q1 = 16'h670e; // 0x1eea
	13'h0f76: q1 = 16'h3ebc; // 0x1eec
	13'h0f77: q1 = 16'h0001; // 0x1eee
	13'h0f78: q1 = 16'h2f0d; // 0x1ef0
	13'h0f79: q1 = 16'h4eb9; // 0x1ef2
	13'h0f7a: q1 = 16'h0000; // 0x1ef4
	13'h0f7b: q1 = 16'h5f04; // 0x1ef6
	13'h0f7c: q1 = 16'h4a9f; // 0x1ef8
	13'h0f7d: q1 = 16'h4a9f; // 0x1efa
	13'h0f7e: q1 = 16'h4cdf; // 0x1efc
	13'h0f7f: q1 = 16'h2080; // 0x1efe
	13'h0f80: q1 = 16'h4e5e; // 0x1f00
	13'h0f81: q1 = 16'h4e75; // 0x1f02
	13'h0f82: q1 = 16'h4e56; // 0x1f04
	13'h0f83: q1 = 16'h0000; // 0x1f06
	13'h0f84: q1 = 16'h48e7; // 0x1f08
	13'h0f85: q1 = 16'h0704; // 0x1f0a
	13'h0f86: q1 = 16'h2a6e; // 0x1f0c
	13'h0f87: q1 = 16'h0008; // 0x1f0e
	13'h0f88: q1 = 16'h3b6e; // 0x1f10
	13'h0f89: q1 = 16'h000c; // 0x1f12
	13'h0f8a: q1 = 16'h0004; // 0x1f14
	13'h0f8b: q1 = 16'h0c6e; // 0x1f16
	13'h0f8c: q1 = 16'h0001; // 0x1f18
	13'h0f8d: q1 = 16'h000c; // 0x1f1a
	13'h0f8e: q1 = 16'h6604; // 0x1f1c
	13'h0f8f: q1 = 16'h7e1e; // 0x1f1e
	13'h0f90: q1 = 16'h6002; // 0x1f20
	13'h0f91: q1 = 16'h7e1c; // 0x1f22
	13'h0f92: q1 = 16'h3c15; // 0x1f24
	13'h0f93: q1 = 16'h3015; // 0x1f26
	13'h0f94: q1 = 16'hd07c; // 0x1f28
	13'h0f95: q1 = 16'h0400; // 0x1f2a
	13'h0f96: q1 = 16'hb046; // 0x1f2c
	13'h0f97: q1 = 16'h6d1c; // 0x1f2e
	13'h0f98: q1 = 16'h3ebc; // 0x1f30
	13'h0f99: q1 = 16'h002a; // 0x1f32
	13'h0f9a: q1 = 16'h3f07; // 0x1f34
	13'h0f9b: q1 = 16'h3f2d; // 0x1f36
	13'h0f9c: q1 = 16'h0002; // 0x1f38
	13'h0f9d: q1 = 16'h3f06; // 0x1f3a
	13'h0f9e: q1 = 16'h4eb9; // 0x1f3c
	13'h0f9f: q1 = 16'h0000; // 0x1f3e
	13'h0fa0: q1 = 16'h3f80; // 0x1f40
	13'h0fa1: q1 = 16'h5c4f; // 0x1f42
	13'h0fa2: q1 = 16'h5247; // 0x1f44
	13'h0fa3: q1 = 16'hdc7c; // 0x1f46
	13'h0fa4: q1 = 16'h0400; // 0x1f48
	13'h0fa5: q1 = 16'h60da; // 0x1f4a
	13'h0fa6: q1 = 16'h4a9f; // 0x1f4c
	13'h0fa7: q1 = 16'h4cdf; // 0x1f4e
	13'h0fa8: q1 = 16'h20c0; // 0x1f50
	13'h0fa9: q1 = 16'h4e5e; // 0x1f52
	13'h0faa: q1 = 16'h4e75; // 0x1f54
	13'h0fab: q1 = 16'h4e56; // 0x1f56
	13'h0fac: q1 = 16'h0000; // 0x1f58
	13'h0fad: q1 = 16'h48e7; // 0x1f5a
	13'h0fae: q1 = 16'h011c; // 0x1f5c
	13'h0faf: q1 = 16'h2a6e; // 0x1f5e
	13'h0fb0: q1 = 16'h0008; // 0x1f60
	13'h0fb1: q1 = 16'h286e; // 0x1f62
	13'h0fb2: q1 = 16'h000c; // 0x1f64
	13'h0fb3: q1 = 16'h266e; // 0x1f66
	13'h0fb4: q1 = 16'h0010; // 0x1f68
	13'h0fb5: q1 = 16'h4a79; // 0x1f6a
	13'h0fb6: q1 = 16'h0001; // 0x1f6c
	13'h0fb7: q1 = 16'h8676; // 0x1f6e
	13'h0fb8: q1 = 16'h666e; // 0x1f70
	13'h0fb9: q1 = 16'h4a79; // 0x1f72
	13'h0fba: q1 = 16'h0001; // 0x1f74
	13'h0fbb: q1 = 16'h7faa; // 0x1f76
	13'h0fbc: q1 = 16'h6666; // 0x1f78
	13'h0fbd: q1 = 16'h2039; // 0x1f7a
	13'h0fbe: q1 = 16'h0001; // 0x1f7c
	13'h0fbf: q1 = 16'h86ae; // 0x1f7e
	13'h0fc0: q1 = 16'h2040; // 0x1f80
	13'h0fc1: q1 = 16'h3215; // 0x1f82
	13'h0fc2: q1 = 16'hc27c; // 0x1f84
	13'h0fc3: q1 = 16'h007f; // 0x1f86
	13'h0fc4: q1 = 16'h1081; // 0x1f88
	13'h0fc5: q1 = 16'h4a54; // 0x1f8a
	13'h0fc6: q1 = 16'h6712; // 0x1f8c
	13'h0fc7: q1 = 16'h3f3c; // 0x1f8e
	13'h0fc8: q1 = 16'h0080; // 0x1f90
	13'h0fc9: q1 = 16'h2039; // 0x1f92
	13'h0fca: q1 = 16'h0001; // 0x1f94
	13'h0fcb: q1 = 16'h86ae; // 0x1f96
	13'h0fcc: q1 = 16'h2040; // 0x1f98
	13'h0fcd: q1 = 16'h1210; // 0x1f9a
	13'h0fce: q1 = 16'h825f; // 0x1f9c
	13'h0fcf: q1 = 16'h1081; // 0x1f9e
	13'h0fd0: q1 = 16'h7001; // 0x1fa0
	13'h0fd1: q1 = 16'h4281; // 0x1fa2
	13'h0fd2: q1 = 16'h3239; // 0x1fa4
	13'h0fd3: q1 = 16'h0001; // 0x1fa6
	13'h0fd4: q1 = 16'h7ba2; // 0x1fa8
	13'h0fd5: q1 = 16'he360; // 0x1faa
	13'h0fd6: q1 = 16'h4640; // 0x1fac
	13'h0fd7: q1 = 16'h3f00; // 0x1fae
	13'h0fd8: q1 = 16'h2039; // 0x1fb0
	13'h0fd9: q1 = 16'h0001; // 0x1fb2
	13'h0fda: q1 = 16'h7ebc; // 0x1fb4
	13'h0fdb: q1 = 16'h2040; // 0x1fb6
	13'h0fdc: q1 = 16'h1210; // 0x1fb8
	13'h0fdd: q1 = 16'hc25f; // 0x1fba
	13'h0fde: q1 = 16'h1081; // 0x1fbc
	13'h0fdf: q1 = 16'h4a53; // 0x1fbe
	13'h0fe0: q1 = 16'h671c; // 0x1fc0
	13'h0fe1: q1 = 16'h7001; // 0x1fc2
	13'h0fe2: q1 = 16'h4281; // 0x1fc4
	13'h0fe3: q1 = 16'h3239; // 0x1fc6
	13'h0fe4: q1 = 16'h0001; // 0x1fc8
	13'h0fe5: q1 = 16'h7ba2; // 0x1fca
	13'h0fe6: q1 = 16'he360; // 0x1fcc
	13'h0fe7: q1 = 16'h3f00; // 0x1fce
	13'h0fe8: q1 = 16'h2039; // 0x1fd0
	13'h0fe9: q1 = 16'h0001; // 0x1fd2
	13'h0fea: q1 = 16'h7ebc; // 0x1fd4
	13'h0feb: q1 = 16'h2040; // 0x1fd6
	13'h0fec: q1 = 16'h1210; // 0x1fd8
	13'h0fed: q1 = 16'h825f; // 0x1fda
	13'h0fee: q1 = 16'h1081; // 0x1fdc
	13'h0fef: q1 = 16'h6050; // 0x1fde
	13'h0ff0: q1 = 16'h2039; // 0x1fe0
	13'h0ff1: q1 = 16'h0001; // 0x1fe2
	13'h0ff2: q1 = 16'h86ae; // 0x1fe4
	13'h0ff3: q1 = 16'h2040; // 0x1fe6
	13'h0ff4: q1 = 16'h1010; // 0x1fe8
	13'h0ff5: q1 = 16'h4880; // 0x1fea
	13'h0ff6: q1 = 16'hc07c; // 0x1fec
	13'h0ff7: q1 = 16'h007f; // 0x1fee
	13'h0ff8: q1 = 16'h3a80; // 0x1ff0
	13'h0ff9: q1 = 16'h2039; // 0x1ff2
	13'h0ffa: q1 = 16'h0001; // 0x1ff4
	13'h0ffb: q1 = 16'h86ae; // 0x1ff6
	13'h0ffc: q1 = 16'h2040; // 0x1ff8
	13'h0ffd: q1 = 16'h1010; // 0x1ffa
	13'h0ffe: q1 = 16'h4880; // 0x1ffc
	13'h0fff: q1 = 16'hc07c; // 0x1ffe
	13'h1000: q1 = 16'h0080; // 0x2000
	13'h1001: q1 = 16'h6604; // 0x2002
	13'h1002: q1 = 16'h4254; // 0x2004
	13'h1003: q1 = 16'h6004; // 0x2006
	13'h1004: q1 = 16'h38bc; // 0x2008
	13'h1005: q1 = 16'h0001; // 0x200a
	13'h1006: q1 = 16'h2039; // 0x200c
	13'h1007: q1 = 16'h0001; // 0x200e
	13'h1008: q1 = 16'h7ebc; // 0x2010
	13'h1009: q1 = 16'h2040; // 0x2012
	13'h100a: q1 = 16'h1010; // 0x2014
	13'h100b: q1 = 16'h4880; // 0x2016
	13'h100c: q1 = 16'h4281; // 0x2018
	13'h100d: q1 = 16'h3239; // 0x201a
	13'h100e: q1 = 16'h0001; // 0x201c
	13'h100f: q1 = 16'h7ba2; // 0x201e
	13'h1010: q1 = 16'he260; // 0x2020
	13'h1011: q1 = 16'hc07c; // 0x2022
	13'h1012: q1 = 16'h0001; // 0x2024
	13'h1013: q1 = 16'h6604; // 0x2026
	13'h1014: q1 = 16'h4253; // 0x2028
	13'h1015: q1 = 16'h6004; // 0x202a
	13'h1016: q1 = 16'h36bc; // 0x202c
	13'h1017: q1 = 16'h0001; // 0x202e
	13'h1018: q1 = 16'h4a79; // 0x2030
	13'h1019: q1 = 16'h0001; // 0x2032
	13'h101a: q1 = 16'h7faa; // 0x2034
	13'h101b: q1 = 16'h6716; // 0x2036
	13'h101c: q1 = 16'h7001; // 0x2038
	13'h101d: q1 = 16'h9079; // 0x203a
	13'h101e: q1 = 16'h0001; // 0x203c
	13'h101f: q1 = 16'h7ba4; // 0x203e
	13'h1020: q1 = 16'h33c0; // 0x2040
	13'h1021: q1 = 16'h0001; // 0x2042
	13'h1022: q1 = 16'h7ba4; // 0x2044
	13'h1023: q1 = 16'h4a79; // 0x2046
	13'h1024: q1 = 16'h0001; // 0x2048
	13'h1025: q1 = 16'h7ba4; // 0x204a
	13'h1026: q1 = 16'h6622; // 0x204c
	13'h1027: q1 = 16'h52b9; // 0x204e
	13'h1028: q1 = 16'h0001; // 0x2050
	13'h1029: q1 = 16'h86ae; // 0x2052
	13'h102a: q1 = 16'h5279; // 0x2054
	13'h102b: q1 = 16'h0001; // 0x2056
	13'h102c: q1 = 16'h7ba2; // 0x2058
	13'h102d: q1 = 16'h0c79; // 0x205a
	13'h102e: q1 = 16'h0007; // 0x205c
	13'h102f: q1 = 16'h0001; // 0x205e
	13'h1030: q1 = 16'h7ba2; // 0x2060
	13'h1031: q1 = 16'h6f0c; // 0x2062
	13'h1032: q1 = 16'h4279; // 0x2064
	13'h1033: q1 = 16'h0001; // 0x2066
	13'h1034: q1 = 16'h7ba2; // 0x2068
	13'h1035: q1 = 16'h52b9; // 0x206a
	13'h1036: q1 = 16'h0001; // 0x206c
	13'h1037: q1 = 16'h7ebc; // 0x206e
	13'h1038: q1 = 16'h4a9f; // 0x2070
	13'h1039: q1 = 16'h4cdf; // 0x2072
	13'h103a: q1 = 16'h3800; // 0x2074
	13'h103b: q1 = 16'h4e5e; // 0x2076
	13'h103c: q1 = 16'h4e75; // 0x2078
	13'h103d: q1 = 16'h4e56; // 0x207a
	13'h103e: q1 = 16'hfffc; // 0x207c
	13'h103f: q1 = 16'h48e7; // 0x207e
	13'h1040: q1 = 16'h3f04; // 0x2080
	13'h1041: q1 = 16'h2a7c; // 0x2082
	13'h1042: q1 = 16'h0001; // 0x2084
	13'h1043: q1 = 16'h7f2c; // 0x2086
	13'h1044: q1 = 16'h4aad; // 0x2088
	13'h1045: q1 = 16'h0006; // 0x208a
	13'h1046: q1 = 16'h6628; // 0x208c
	13'h1047: q1 = 16'h4aad; // 0x208e
	13'h1048: q1 = 16'h001c; // 0x2090
	13'h1049: q1 = 16'h6622; // 0x2092
	13'h104a: q1 = 16'h4245; // 0x2094
	13'h104b: q1 = 16'h4a6d; // 0x2096
	13'h104c: q1 = 16'h0010; // 0x2098
	13'h104d: q1 = 16'h6712; // 0x209a
	13'h104e: q1 = 16'h3015; // 0x209c
	13'h104f: q1 = 16'h48c0; // 0x209e
	13'h1050: q1 = 16'hd0bc; // 0x20a0
	13'h1051: q1 = 16'h0000; // 0x20a2
	13'h1052: q1 = 16'hcb52; // 0x20a4
	13'h1053: q1 = 16'h2040; // 0x20a6
	13'h1054: q1 = 16'h1e10; // 0x20a8
	13'h1055: q1 = 16'h4887; // 0x20aa
	13'h1056: q1 = 16'h6004; // 0x20ac
	13'h1057: q1 = 16'h3e3c; // 0x20ae
	13'h1058: q1 = 16'h00be; // 0x20b0
	13'h1059: q1 = 16'h6000; // 0x20b2
	13'h105a: q1 = 16'h00f8; // 0x20b4
	13'h105b: q1 = 16'h4aad; // 0x20b6
	13'h105c: q1 = 16'h001c; // 0x20b8
	13'h105d: q1 = 16'h6f38; // 0x20ba
	13'h105e: q1 = 16'h0cad; // 0x20bc
	13'h105f: q1 = 16'h0000; // 0x20be
	13'h1060: q1 = 16'h0005; // 0x20c0
	13'h1061: q1 = 16'h001c; // 0x20c2
	13'h1062: q1 = 16'h6c2e; // 0x20c4
	13'h1063: q1 = 16'h2039; // 0x20c6
	13'h1064: q1 = 16'h0000; // 0x20c8
	13'h1065: q1 = 16'hcc5a; // 0x20ca
	13'h1066: q1 = 16'h90ad; // 0x20cc
	13'h1067: q1 = 16'h001c; // 0x20ce
	13'h1068: q1 = 16'h3e00; // 0x20d0
	13'h1069: q1 = 16'hde7c; // 0x20d2
	13'h106a: q1 = 16'h0050; // 0x20d4
	13'h106b: q1 = 16'h3a3c; // 0x20d6
	13'h106c: q1 = 16'h0080; // 0x20d8
	13'h106d: q1 = 16'h4a79; // 0x20da
	13'h106e: q1 = 16'h0001; // 0x20dc
	13'h106f: q1 = 16'h7f20; // 0x20de
	13'h1070: q1 = 16'h6708; // 0x20e0
	13'h1071: q1 = 16'h4244; // 0x20e2
	13'h1072: q1 = 16'h363c; // 0x20e4
	13'h1073: q1 = 16'h0400; // 0x20e6
	13'h1074: q1 = 16'h6008; // 0x20e8
	13'h1075: q1 = 16'h383c; // 0x20ea
	13'h1076: q1 = 16'hfc00; // 0x20ec
	13'h1077: q1 = 16'h363c; // 0x20ee
	13'h1078: q1 = 16'h0380; // 0x20f0
	13'h1079: q1 = 16'h6058; // 0x20f2
	13'h107a: q1 = 16'h302d; // 0x20f4
	13'h107b: q1 = 16'h000e; // 0x20f6
	13'h107c: q1 = 16'h48c0; // 0x20f8
	13'h107d: q1 = 16'hd0bc; // 0x20fa
	13'h107e: q1 = 16'h0000; // 0x20fc
	13'h107f: q1 = 16'hca18; // 0x20fe
	13'h1080: q1 = 16'h2040; // 0x2100
	13'h1081: q1 = 16'h1e10; // 0x2102
	13'h1082: q1 = 16'h4887; // 0x2104
	13'h1083: q1 = 16'hde7c; // 0x2106
	13'h1084: q1 = 16'h00ec; // 0x2108
	13'h1085: q1 = 16'h3c07; // 0x210a
	13'h1086: q1 = 16'hdc7c; // 0x210c
	13'h1087: q1 = 16'hff14; // 0x210e
	13'h1088: q1 = 16'h3006; // 0x2110
	13'h1089: q1 = 16'h48c0; // 0x2112
	13'h108a: q1 = 16'hd0bc; // 0x2114
	13'h108b: q1 = 16'h0000; // 0x2116
	13'h108c: q1 = 16'hcc4c; // 0x2118
	13'h108d: q1 = 16'h2040; // 0x211a
	13'h108e: q1 = 16'h1a10; // 0x211c
	13'h108f: q1 = 16'h4885; // 0x211e
	13'h1090: q1 = 16'hef45; // 0x2120
	13'h1091: q1 = 16'h3006; // 0x2122
	13'h1092: q1 = 16'h48c0; // 0x2124
	13'h1093: q1 = 16'hd0bc; // 0x2126
	13'h1094: q1 = 16'h0000; // 0x2128
	13'h1095: q1 = 16'hcc30; // 0x212a
	13'h1096: q1 = 16'h2040; // 0x212c
	13'h1097: q1 = 16'h1810; // 0x212e
	13'h1098: q1 = 16'h4884; // 0x2130
	13'h1099: q1 = 16'hef44; // 0x2132
	13'h109a: q1 = 16'h3004; // 0x2134
	13'h109b: q1 = 16'h4440; // 0x2136
	13'h109c: q1 = 16'h3800; // 0x2138
	13'h109d: q1 = 16'h3006; // 0x213a
	13'h109e: q1 = 16'h48c0; // 0x213c
	13'h109f: q1 = 16'hd0bc; // 0x213e
	13'h10a0: q1 = 16'h0000; // 0x2140
	13'h10a1: q1 = 16'hcc3e; // 0x2142
	13'h10a2: q1 = 16'h2040; // 0x2144
	13'h10a3: q1 = 16'h1610; // 0x2146
	13'h10a4: q1 = 16'h4883; // 0x2148
	13'h10a5: q1 = 16'hef43; // 0x214a
	13'h10a6: q1 = 16'h0c6d; // 0x214c
	13'h10a7: q1 = 16'h0012; // 0x214e
	13'h10a8: q1 = 16'h000e; // 0x2150
	13'h10a9: q1 = 16'h6f14; // 0x2152
	13'h10aa: q1 = 16'h0c6d; // 0x2154
	13'h10ab: q1 = 16'h0036; // 0x2156
	13'h10ac: q1 = 16'h000e; // 0x2158
	13'h10ad: q1 = 16'h6e0c; // 0x215a
	13'h10ae: q1 = 16'h3005; // 0x215c
	13'h10af: q1 = 16'h4440; // 0x215e
	13'h10b0: q1 = 16'h3a00; // 0x2160
	13'h10b1: q1 = 16'h3004; // 0x2162
	13'h10b2: q1 = 16'h4440; // 0x2164
	13'h10b3: q1 = 16'h3800; // 0x2166
	13'h10b4: q1 = 16'h4aad; // 0x2168
	13'h10b5: q1 = 16'h0006; // 0x216a
	13'h10b6: q1 = 16'h673e; // 0x216c
	13'h10b7: q1 = 16'h206d; // 0x216e
	13'h10b8: q1 = 16'h0024; // 0x2170
	13'h10b9: q1 = 16'h3010; // 0x2172
	13'h10ba: q1 = 16'hd044; // 0x2174
	13'h10bb: q1 = 16'h3d40; // 0x2176
	13'h10bc: q1 = 16'hfffe; // 0x2178
	13'h10bd: q1 = 16'h206d; // 0x217a
	13'h10be: q1 = 16'h0024; // 0x217c
	13'h10bf: q1 = 16'h3028; // 0x217e
	13'h10c0: q1 = 16'h0002; // 0x2180
	13'h10c1: q1 = 16'hd043; // 0x2182
	13'h10c2: q1 = 16'h3d40; // 0x2184
	13'h10c3: q1 = 16'hfffc; // 0x2186
	13'h10c4: q1 = 16'h202d; // 0x2188
	13'h10c5: q1 = 16'h001c; // 0x218a
	13'h10c6: q1 = 16'h4a40; // 0x218c
	13'h10c7: q1 = 16'h6704; // 0x218e
	13'h10c8: q1 = 16'h4257; // 0x2190
	13'h10c9: q1 = 16'h6004; // 0x2192
	13'h10ca: q1 = 16'h3ebc; // 0x2194
	13'h10cb: q1 = 16'h0001; // 0x2196
	13'h10cc: q1 = 16'h3f2e; // 0x2198
	13'h10cd: q1 = 16'hfffc; // 0x219a
	13'h10ce: q1 = 16'h3f2e; // 0x219c
	13'h10cf: q1 = 16'hfffe; // 0x219e
	13'h10d0: q1 = 16'h2f2d; // 0x21a0
	13'h10d1: q1 = 16'h0006; // 0x21a2
	13'h10d2: q1 = 16'h4eb9; // 0x21a4
	13'h10d3: q1 = 16'h0000; // 0x21a6
	13'h10d4: q1 = 16'h3c92; // 0x21a8
	13'h10d5: q1 = 16'hbf8f; // 0x21aa
	13'h10d6: q1 = 16'h206d; // 0x21ac
	13'h10d7: q1 = 16'h0028; // 0x21ae
	13'h10d8: q1 = 16'h226d; // 0x21b0
	13'h10d9: q1 = 16'h0024; // 0x21b2
	13'h10da: q1 = 16'h3211; // 0x21b4
	13'h10db: q1 = 16'hd245; // 0x21b6
	13'h10dc: q1 = 16'h3081; // 0x21b8
	13'h10dd: q1 = 16'h206d; // 0x21ba
	13'h10de: q1 = 16'h0028; // 0x21bc
	13'h10df: q1 = 16'h226d; // 0x21be
	13'h10e0: q1 = 16'h0024; // 0x21c0
	13'h10e1: q1 = 16'h3169; // 0x21c2
	13'h10e2: q1 = 16'h0002; // 0x21c4
	13'h10e3: q1 = 16'h0002; // 0x21c6
	13'h10e4: q1 = 16'h206d; // 0x21c8
	13'h10e5: q1 = 16'h0028; // 0x21ca
	13'h10e6: q1 = 16'h3147; // 0x21cc
	13'h10e7: q1 = 16'h0004; // 0x21ce
	13'h10e8: q1 = 16'h206d; // 0x21d0
	13'h10e9: q1 = 16'h0028; // 0x21d2
	13'h10ea: q1 = 16'h317c; // 0x21d4
	13'h10eb: q1 = 16'h0015; // 0x21d6
	13'h10ec: q1 = 16'h0006; // 0x21d8
	13'h10ed: q1 = 16'h3ead; // 0x21da
	13'h10ee: q1 = 16'h000e; // 0x21dc
	13'h10ef: q1 = 16'h202d; // 0x21de
	13'h10f0: q1 = 16'h0028; // 0x21e0
	13'h10f1: q1 = 16'h5c80; // 0x21e2
	13'h10f2: q1 = 16'h2f00; // 0x21e4
	13'h10f3: q1 = 16'h4eb9; // 0x21e6
	13'h10f4: q1 = 16'h0000; // 0x21e8
	13'h10f5: q1 = 16'h3ee6; // 0x21ea
	13'h10f6: q1 = 16'h4a9f; // 0x21ec
	13'h10f7: q1 = 16'h4a9f; // 0x21ee
	13'h10f8: q1 = 16'h4cdf; // 0x21f0
	13'h10f9: q1 = 16'h20f8; // 0x21f2
	13'h10fa: q1 = 16'h4e5e; // 0x21f4
	13'h10fb: q1 = 16'h4e75; // 0x21f6
	13'h10fc: q1 = 16'h4e56; // 0x21f8
	13'h10fd: q1 = 16'h0000; // 0x21fa
	13'h10fe: q1 = 16'h48e7; // 0x21fc
	13'h10ff: q1 = 16'h0304; // 0x21fe
	13'h1100: q1 = 16'h2a7c; // 0x2200
	13'h1101: q1 = 16'h0001; // 0x2202
	13'h1102: q1 = 16'h7f2c; // 0x2204
	13'h1103: q1 = 16'h206d; // 0x2206
	13'h1104: q1 = 16'h0024; // 0x2208
	13'h1105: q1 = 16'h3b68; // 0x220a
	13'h1106: q1 = 16'h0002; // 0x220c
	13'h1107: q1 = 16'h0030; // 0x220e
	13'h1108: q1 = 16'h206d; // 0x2210
	13'h1109: q1 = 16'h0020; // 0x2212
	13'h110a: q1 = 16'h226d; // 0x2214
	13'h110b: q1 = 16'h0024; // 0x2216
	13'h110c: q1 = 16'h3091; // 0x2218
	13'h110d: q1 = 16'h206d; // 0x221a
	13'h110e: q1 = 16'h002c; // 0x221c
	13'h110f: q1 = 16'h226d; // 0x221e
	13'h1110: q1 = 16'h0020; // 0x2220
	13'h1111: q1 = 16'h3091; // 0x2222
	13'h1112: q1 = 16'h206d; // 0x2224
	13'h1113: q1 = 16'h0020; // 0x2226
	13'h1114: q1 = 16'h226d; // 0x2228
	13'h1115: q1 = 16'h0024; // 0x222a
	13'h1116: q1 = 16'h3229; // 0x222c
	13'h1117: q1 = 16'h0002; // 0x222e
	13'h1118: q1 = 16'hd27c; // 0x2230
	13'h1119: q1 = 16'h0200; // 0x2232
	13'h111a: q1 = 16'h3141; // 0x2234
	13'h111b: q1 = 16'h0002; // 0x2236
	13'h111c: q1 = 16'h206d; // 0x2238
	13'h111d: q1 = 16'h002c; // 0x223a
	13'h111e: q1 = 16'h226d; // 0x223c
	13'h111f: q1 = 16'h0020; // 0x223e
	13'h1120: q1 = 16'h3169; // 0x2240
	13'h1121: q1 = 16'h0002; // 0x2242
	13'h1122: q1 = 16'h0002; // 0x2244
	13'h1123: q1 = 16'h206d; // 0x2246
	13'h1124: q1 = 16'h0024; // 0x2248
	13'h1125: q1 = 16'h317c; // 0x224a
	13'h1126: q1 = 16'h0005; // 0x224c
	13'h1127: q1 = 16'h0006; // 0x224e
	13'h1128: q1 = 16'h206d; // 0x2250
	13'h1129: q1 = 16'h0020; // 0x2252
	13'h112a: q1 = 16'h317c; // 0x2254
	13'h112b: q1 = 16'h0007; // 0x2256
	13'h112c: q1 = 16'h0006; // 0x2258
	13'h112d: q1 = 16'h206d; // 0x225a
	13'h112e: q1 = 16'h002c; // 0x225c
	13'h112f: q1 = 16'h317c; // 0x225e
	13'h1130: q1 = 16'h001d; // 0x2260
	13'h1131: q1 = 16'h0006; // 0x2262
	13'h1132: q1 = 16'h4255; // 0x2264
	13'h1133: q1 = 16'h426d; // 0x2266
	13'h1134: q1 = 16'h0012; // 0x2268
	13'h1135: q1 = 16'h426d; // 0x226a
	13'h1136: q1 = 16'h0018; // 0x226c
	13'h1137: q1 = 16'h426d; // 0x226e
	13'h1138: q1 = 16'h001a; // 0x2270
	13'h1139: q1 = 16'h42ad; // 0x2272
	13'h113a: q1 = 16'h001c; // 0x2274
	13'h113b: q1 = 16'h426d; // 0x2276
	13'h113c: q1 = 16'h0010; // 0x2278
	13'h113d: q1 = 16'h3b7c; // 0x227a
	13'h113e: q1 = 16'h0002; // 0x227c
	13'h113f: q1 = 16'h0004; // 0x227e
	13'h1140: q1 = 16'h3b6d; // 0x2280
	13'h1141: q1 = 16'h0004; // 0x2282
	13'h1142: q1 = 16'h0002; // 0x2284
	13'h1143: q1 = 16'h2b79; // 0x2286
	13'h1144: q1 = 16'h0000; // 0x2288
	13'h1145: q1 = 16'hcc5e; // 0x228a
	13'h1146: q1 = 16'h000a; // 0x228c
	13'h1147: q1 = 16'h206d; // 0x228e
	13'h1148: q1 = 16'h0024; // 0x2290
	13'h1149: q1 = 16'h317c; // 0x2292
	13'h114a: q1 = 16'h00bf; // 0x2294
	13'h114b: q1 = 16'h0004; // 0x2296
	13'h114c: q1 = 16'h3ead; // 0x2298
	13'h114d: q1 = 16'h000e; // 0x229a
	13'h114e: q1 = 16'h202d; // 0x229c
	13'h114f: q1 = 16'h0024; // 0x229e
	13'h1150: q1 = 16'h5c80; // 0x22a0
	13'h1151: q1 = 16'h2f00; // 0x22a2
	13'h1152: q1 = 16'h4eb9; // 0x22a4
	13'h1153: q1 = 16'h0000; // 0x22a6
	13'h1154: q1 = 16'h3ee6; // 0x22a8
	13'h1155: q1 = 16'h4a9f; // 0x22aa
	13'h1156: q1 = 16'h302d; // 0x22ac
	13'h1157: q1 = 16'h000e; // 0x22ae
	13'h1158: q1 = 16'h48c0; // 0x22b0
	13'h1159: q1 = 16'hd0bc; // 0x22b2
	13'h115a: q1 = 16'h0000; // 0x22b4
	13'h115b: q1 = 16'hca18; // 0x22b6
	13'h115c: q1 = 16'h2040; // 0x22b8
	13'h115d: q1 = 16'h1e10; // 0x22ba
	13'h115e: q1 = 16'h4887; // 0x22bc
	13'h115f: q1 = 16'h206d; // 0x22be
	13'h1160: q1 = 16'h0020; // 0x22c0
	13'h1161: q1 = 16'h3207; // 0x22c2
	13'h1162: q1 = 16'hd27c; // 0x22c4
	13'h1163: q1 = 16'h000c; // 0x22c6
	13'h1164: q1 = 16'h3141; // 0x22c8
	13'h1165: q1 = 16'h0004; // 0x22ca
	13'h1166: q1 = 16'h3ead; // 0x22cc
	13'h1167: q1 = 16'h000e; // 0x22ce
	13'h1168: q1 = 16'h202d; // 0x22d0
	13'h1169: q1 = 16'h0020; // 0x22d2
	13'h116a: q1 = 16'h5c80; // 0x22d4
	13'h116b: q1 = 16'h2f00; // 0x22d6
	13'h116c: q1 = 16'h4eb9; // 0x22d8
	13'h116d: q1 = 16'h0000; // 0x22da
	13'h116e: q1 = 16'h3ee6; // 0x22dc
	13'h116f: q1 = 16'h4a9f; // 0x22de
	13'h1170: q1 = 16'h206d; // 0x22e0
	13'h1171: q1 = 16'h002c; // 0x22e2
	13'h1172: q1 = 16'h3207; // 0x22e4
	13'h1173: q1 = 16'h48c1; // 0x22e6
	13'h1174: q1 = 16'hd2bc; // 0x22e8
	13'h1175: q1 = 16'h0000; // 0x22ea
	13'h1176: q1 = 16'hcb62; // 0x22ec
	13'h1177: q1 = 16'h2241; // 0x22ee
	13'h1178: q1 = 16'h1211; // 0x22f0
	13'h1179: q1 = 16'h4881; // 0x22f2
	13'h117a: q1 = 16'h3141; // 0x22f4
	13'h117b: q1 = 16'h0004; // 0x22f6
	13'h117c: q1 = 16'h3ead; // 0x22f8
	13'h117d: q1 = 16'h000e; // 0x22fa
	13'h117e: q1 = 16'h202d; // 0x22fc
	13'h117f: q1 = 16'h002c; // 0x22fe
	13'h1180: q1 = 16'h5c80; // 0x2300
	13'h1181: q1 = 16'h2f00; // 0x2302
	13'h1182: q1 = 16'h4eb9; // 0x2304
	13'h1183: q1 = 16'h0000; // 0x2306
	13'h1184: q1 = 16'h3ee6; // 0x2308
	13'h1185: q1 = 16'h4a9f; // 0x230a
	13'h1186: q1 = 16'h4a9f; // 0x230c
	13'h1187: q1 = 16'h4cdf; // 0x230e
	13'h1188: q1 = 16'h2080; // 0x2310
	13'h1189: q1 = 16'h4e5e; // 0x2312
	13'h118a: q1 = 16'h4e75; // 0x2314
	13'h118b: q1 = 16'h4e56; // 0x2316
	13'h118c: q1 = 16'h0000; // 0x2318
	13'h118d: q1 = 16'h48e7; // 0x231a
	13'h118e: q1 = 16'h031c; // 0x231c
	13'h118f: q1 = 16'h33fc; // 0x231e
	13'h1190: q1 = 16'h002d; // 0x2320
	13'h1191: q1 = 16'h0001; // 0x2322
	13'h1192: q1 = 16'h893c; // 0x2324
	13'h1193: q1 = 16'h4eb9; // 0x2326
	13'h1194: q1 = 16'h0000; // 0x2328
	13'h1195: q1 = 16'h01de; // 0x232a
	13'h1196: q1 = 16'h4279; // 0x232c
	13'h1197: q1 = 16'h0001; // 0x232e
	13'h1198: q1 = 16'h8a7c; // 0x2330
	13'h1199: q1 = 16'h42b9; // 0x2332
	13'h119a: q1 = 16'h0001; // 0x2334
	13'h119b: q1 = 16'h7f60; // 0x2336
	13'h119c: q1 = 16'h33fc; // 0x2338
	13'h119d: q1 = 16'h0001; // 0x233a
	13'h119e: q1 = 16'h0001; // 0x233c
	13'h119f: q1 = 16'h87dc; // 0x233e
	13'h11a0: q1 = 16'h42b9; // 0x2340
	13'h11a1: q1 = 16'h0001; // 0x2342
	13'h11a2: q1 = 16'h7fac; // 0x2344
	13'h11a3: q1 = 16'h33fc; // 0x2346
	13'h11a4: q1 = 16'h003c; // 0x2348
	13'h11a5: q1 = 16'h0001; // 0x234a
	13'h11a6: q1 = 16'h7fb0; // 0x234c
	13'h11a7: q1 = 16'h42b9; // 0x234e
	13'h11a8: q1 = 16'h0001; // 0x2350
	13'h11a9: q1 = 16'h7fa2; // 0x2352
	13'h11aa: q1 = 16'h4279; // 0x2354
	13'h11ab: q1 = 16'h0001; // 0x2356
	13'h11ac: q1 = 16'h7590; // 0x2358
	13'h11ad: q1 = 16'h42b9; // 0x235a
	13'h11ae: q1 = 16'h0001; // 0x235c
	13'h11af: q1 = 16'h7fc2; // 0x235e
	13'h11b0: q1 = 16'h33fc; // 0x2360
	13'h11b1: q1 = 16'h7400; // 0x2362
	13'h11b2: q1 = 16'h0001; // 0x2364
	13'h11b3: q1 = 16'h8662; // 0x2366
	13'h11b4: q1 = 16'h33fc; // 0x2368
	13'h11b5: q1 = 16'h7c00; // 0x236a
	13'h11b6: q1 = 16'h0001; // 0x236c
	13'h11b7: q1 = 16'h8664; // 0x236e
	13'h11b8: q1 = 16'h33fc; // 0x2370
	13'h11b9: q1 = 16'h7c00; // 0x2372
	13'h11ba: q1 = 16'h0001; // 0x2374
	13'h11bb: q1 = 16'h863e; // 0x2376
	13'h11bc: q1 = 16'h4eb9; // 0x2378
	13'h11bd: q1 = 16'h0000; // 0x237a
	13'h11be: q1 = 16'h0226; // 0x237c
	13'h11bf: q1 = 16'h4279; // 0x237e
	13'h11c0: q1 = 16'h0001; // 0x2380
	13'h11c1: q1 = 16'h7f5e; // 0x2382
	13'h11c2: q1 = 16'h4279; // 0x2384
	13'h11c3: q1 = 16'h0001; // 0x2386
	13'h11c4: q1 = 16'h8a7a; // 0x2388
	13'h11c5: q1 = 16'h4279; // 0x238a
	13'h11c6: q1 = 16'h0001; // 0x238c
	13'h11c7: q1 = 16'h7fa6; // 0x238e
	13'h11c8: q1 = 16'h4279; // 0x2390
	13'h11c9: q1 = 16'h0001; // 0x2392
	13'h11ca: q1 = 16'h8052; // 0x2394
	13'h11cb: q1 = 16'h4279; // 0x2396
	13'h11cc: q1 = 16'h0001; // 0x2398
	13'h11cd: q1 = 16'h8676; // 0x239a
	13'h11ce: q1 = 16'h4279; // 0x239c
	13'h11cf: q1 = 16'h0001; // 0x239e
	13'h11d0: q1 = 16'h77e8; // 0x23a0
	13'h11d1: q1 = 16'h33fc; // 0x23a2
	13'h11d2: q1 = 16'h0001; // 0x23a4
	13'h11d3: q1 = 16'h0001; // 0x23a6
	13'h11d4: q1 = 16'h7fc6; // 0x23a8
	13'h11d5: q1 = 16'h4279; // 0x23aa
	13'h11d6: q1 = 16'h0001; // 0x23ac
	13'h11d7: q1 = 16'h7faa; // 0x23ae
	13'h11d8: q1 = 16'h4279; // 0x23b0
	13'h11d9: q1 = 16'h0001; // 0x23b2
	13'h11da: q1 = 16'h806e; // 0x23b4
	13'h11db: q1 = 16'h4279; // 0x23b6
	13'h11dc: q1 = 16'h0001; // 0x23b8
	13'h11dd: q1 = 16'h7bd6; // 0x23ba
	13'h11de: q1 = 16'h4279; // 0x23bc
	13'h11df: q1 = 16'h0001; // 0x23be
	13'h11e0: q1 = 16'h7f2a; // 0x23c0
	13'h11e1: q1 = 16'h4279; // 0x23c2
	13'h11e2: q1 = 16'h0001; // 0x23c4
	13'h11e3: q1 = 16'h7f20; // 0x23c6
	13'h11e4: q1 = 16'h4279; // 0x23c8
	13'h11e5: q1 = 16'h0001; // 0x23ca
	13'h11e6: q1 = 16'h7fa8; // 0x23cc
	13'h11e7: q1 = 16'h23f9; // 0x23ce
	13'h11e8: q1 = 16'h0000; // 0x23d0
	13'h11e9: q1 = 16'hcc62; // 0x23d2
	13'h11ea: q1 = 16'h0001; // 0x23d4
	13'h11eb: q1 = 16'h862c; // 0x23d6
	13'h11ec: q1 = 16'h2ebc; // 0x23d8
	13'h11ed: q1 = 16'h0000; // 0x23da
	13'h11ee: q1 = 16'hcc66; // 0x23dc
	13'h11ef: q1 = 16'h2f3c; // 0x23de
	13'h11f0: q1 = 16'h0001; // 0x23e0
	13'h11f1: q1 = 16'h8630; // 0x23e2
	13'h11f2: q1 = 16'h4eb9; // 0x23e4
	13'h11f3: q1 = 16'h0000; // 0x23e6
	13'h11f4: q1 = 16'h0750; // 0x23e8
	13'h11f5: q1 = 16'h4a9f; // 0x23ea
	13'h11f6: q1 = 16'h267c; // 0x23ec
	13'h11f7: q1 = 16'h0001; // 0x23ee
	13'h11f8: q1 = 16'h8072; // 0x23f0
	13'h11f9: q1 = 16'h4247; // 0x23f2
	13'h11fa: q1 = 16'h2a7c; // 0x23f4
	13'h11fb: q1 = 16'h0001; // 0x23f6
	13'h11fc: q1 = 16'h89be; // 0x23f8
	13'h11fd: q1 = 16'hbe7c; // 0x23fa
	13'h11fe: q1 = 16'h0004; // 0x23fc
	13'h11ff: q1 = 16'h6c44; // 0x23fe
	13'h1200: q1 = 16'h3007; // 0x2400
	13'h1201: q1 = 16'he740; // 0x2402
	13'h1202: q1 = 16'h48c0; // 0x2404
	13'h1203: q1 = 16'hd08b; // 0x2406
	13'h1204: q1 = 16'hd0bc; // 0x2408
	13'h1205: q1 = 16'h0000; // 0x240a
	13'h1206: q1 = 16'h0040; // 0x240c
	13'h1207: q1 = 16'h2b40; // 0x240e
	13'h1208: q1 = 16'h001e; // 0x2410
	13'h1209: q1 = 16'h3007; // 0x2412
	13'h120a: q1 = 16'he740; // 0x2414
	13'h120b: q1 = 16'h48c0; // 0x2416
	13'h120c: q1 = 16'hd08b; // 0x2418
	13'h120d: q1 = 16'hd0bc; // 0x241a
	13'h120e: q1 = 16'h0000; // 0x241c
	13'h120f: q1 = 16'h0060; // 0x241e
	13'h1210: q1 = 16'h2b40; // 0x2420
	13'h1211: q1 = 16'h0022; // 0x2422
	13'h1212: q1 = 16'h3007; // 0x2424
	13'h1213: q1 = 16'he740; // 0x2426
	13'h1214: q1 = 16'h48c0; // 0x2428
	13'h1215: q1 = 16'hd08b; // 0x242a
	13'h1216: q1 = 16'hd0bc; // 0x242c
	13'h1217: q1 = 16'h0000; // 0x242e
	13'h1218: q1 = 16'h0080; // 0x2430
	13'h1219: q1 = 16'h2b40; // 0x2432
	13'h121a: q1 = 16'h0026; // 0x2434
	13'h121b: q1 = 16'h42ad; // 0x2436
	13'h121c: q1 = 16'h0010; // 0x2438
	13'h121d: q1 = 16'h5247; // 0x243a
	13'h121e: q1 = 16'hdbfc; // 0x243c
	13'h121f: q1 = 16'h0000; // 0x243e
	13'h1220: q1 = 16'h002e; // 0x2440
	13'h1221: q1 = 16'h60b6; // 0x2442
	13'h1222: q1 = 16'h41d3; // 0x2444
	13'h1223: q1 = 16'h23c8; // 0x2446
	13'h1224: q1 = 16'h0001; // 0x2448
	13'h1225: q1 = 16'h7f50; // 0x244a
	13'h1226: q1 = 16'h41eb; // 0x244c
	13'h1227: q1 = 16'h0008; // 0x244e
	13'h1228: q1 = 16'h23c8; // 0x2450
	13'h1229: q1 = 16'h0001; // 0x2452
	13'h122a: q1 = 16'h7f4c; // 0x2454
	13'h122b: q1 = 16'h41eb; // 0x2456
	13'h122c: q1 = 16'h0028; // 0x2458
	13'h122d: q1 = 16'h23c8; // 0x245a
	13'h122e: q1 = 16'h0001; // 0x245c
	13'h122f: q1 = 16'h7f54; // 0x245e
	13'h1230: q1 = 16'h41eb; // 0x2460
	13'h1231: q1 = 16'h0030; // 0x2462
	13'h1232: q1 = 16'h23c8; // 0x2464
	13'h1233: q1 = 16'h0001; // 0x2466
	13'h1234: q1 = 16'h7f58; // 0x2468
	13'h1235: q1 = 16'h42b9; // 0x246a
	13'h1236: q1 = 16'h0001; // 0x246c
	13'h1237: q1 = 16'h7f32; // 0x246e
	13'h1238: q1 = 16'h42b9; // 0x2470
	13'h1239: q1 = 16'h0001; // 0x2472
	13'h123a: q1 = 16'h7f36; // 0x2474
	13'h123b: q1 = 16'h4247; // 0x2476
	13'h123c: q1 = 16'h287c; // 0x2478
	13'h123d: q1 = 16'h0001; // 0x247a
	13'h123e: q1 = 16'h7bda; // 0x247c
	13'h123f: q1 = 16'hbe7c; // 0x247e
	13'h1240: q1 = 16'h001a; // 0x2480
	13'h1241: q1 = 16'h6c1c; // 0x2482
	13'h1242: q1 = 16'h3007; // 0x2484
	13'h1243: q1 = 16'he740; // 0x2486
	13'h1244: q1 = 16'h48c0; // 0x2488
	13'h1245: q1 = 16'hd08b; // 0x248a
	13'h1246: q1 = 16'hd0bc; // 0x248c
	13'h1247: q1 = 16'h0000; // 0x248e
	13'h1248: q1 = 16'h00a0; // 0x2490
	13'h1249: q1 = 16'h2940; // 0x2492
	13'h124a: q1 = 16'h0012; // 0x2494
	13'h124b: q1 = 16'h5247; // 0x2496
	13'h124c: q1 = 16'hd9fc; // 0x2498
	13'h124d: q1 = 16'h0000; // 0x249a
	13'h124e: q1 = 16'h001c; // 0x249c
	13'h124f: q1 = 16'h60de; // 0x249e
	13'h1250: q1 = 16'h4eb9; // 0x24a0
	13'h1251: q1 = 16'h0000; // 0x24a2
	13'h1252: q1 = 16'h4754; // 0x24a4
	13'h1253: q1 = 16'h4eb9; // 0x24a6
	13'h1254: q1 = 16'h0000; // 0x24a8
	13'h1255: q1 = 16'h33e6; // 0x24aa
	13'h1256: q1 = 16'h4eb9; // 0x24ac
	13'h1257: q1 = 16'h0000; // 0x24ae
	13'h1258: q1 = 16'h01d8; // 0x24b0
	13'h1259: q1 = 16'h4a9f; // 0x24b2
	13'h125a: q1 = 16'h4cdf; // 0x24b4
	13'h125b: q1 = 16'h3880; // 0x24b6
	13'h125c: q1 = 16'h4e5e; // 0x24b8
	13'h125d: q1 = 16'h4e75; // 0x24ba
	13'h125e: q1 = 16'h4e56; // 0x24bc
	13'h125f: q1 = 16'hffba; // 0x24be
	13'h1260: q1 = 16'h48e7; // 0x24c0
	13'h1261: q1 = 16'h3f04; // 0x24c2
	13'h1262: q1 = 16'h3e2e; // 0x24c4
	13'h1263: q1 = 16'h0008; // 0x24c6
	13'h1264: q1 = 16'h3007; // 0x24c8
	13'h1265: q1 = 16'hc1fc; // 0x24ca
	13'h1266: q1 = 16'h0026; // 0x24cc
	13'h1267: q1 = 16'h2a40; // 0x24ce
	13'h1268: q1 = 16'hdbfc; // 0x24d0
	13'h1269: q1 = 16'h0001; // 0x24d2
	13'h126a: q1 = 16'h8628; // 0x24d4
	13'h126b: q1 = 16'h4a79; // 0x24d6
	13'h126c: q1 = 16'h0001; // 0x24d8
	13'h126d: q1 = 16'h7584; // 0x24da
	13'h126e: q1 = 16'h6738; // 0x24dc
	13'h126f: q1 = 16'h0cad; // 0x24de
	13'h1270: q1 = 16'h0000; // 0x24e0
	13'h1271: q1 = 16'h01f4; // 0x24e2
	13'h1272: q1 = 16'h0004; // 0x24e4
	13'h1273: q1 = 16'h662e; // 0x24e6
	13'h1274: q1 = 16'h2d7c; // 0x24e8
	13'h1275: q1 = 16'h0000; // 0x24ea
	13'h1276: q1 = 16'h0105; // 0x24ec
	13'h1277: q1 = 16'hffba; // 0x24ee
	13'h1278: q1 = 16'h202e; // 0x24f0
	13'h1279: q1 = 16'hffba; // 0x24f2
	13'h127a: q1 = 16'he180; // 0x24f4
	13'h127b: q1 = 16'h2d40; // 0x24f6
	13'h127c: q1 = 16'hffba; // 0x24f8
	13'h127d: q1 = 16'h00ae; // 0x24fa
	13'h127e: q1 = 16'h0000; // 0x24fc
	13'h127f: q1 = 16'h000e; // 0x24fe
	13'h1280: q1 = 16'hffba; // 0x2500
	13'h1281: q1 = 16'h06ae; // 0x2502
	13'h1282: q1 = 16'h0000; // 0x2504
	13'h1283: q1 = 16'h7080; // 0x2506
	13'h1284: q1 = 16'hffba; // 0x2508
	13'h1285: q1 = 16'h202e; // 0x250a
	13'h1286: q1 = 16'hffba; // 0x250c
	13'h1287: q1 = 16'h2040; // 0x250e
	13'h1288: q1 = 16'h117c; // 0x2510
	13'h1289: q1 = 16'h0001; // 0x2512
	13'h128a: q1 = 16'h0001; // 0x2514
	13'h128b: q1 = 16'h4a6d; // 0x2516
	13'h128c: q1 = 16'h001e; // 0x2518
	13'h128d: q1 = 16'h6700; // 0x251a
	13'h128e: q1 = 16'h05a4; // 0x251c
	13'h128f: q1 = 16'h4eb9; // 0x251e
	13'h1290: q1 = 16'h0000; // 0x2520
	13'h1291: q1 = 16'h0226; // 0x2522
	13'h1292: q1 = 16'h4a79; // 0x2524
	13'h1293: q1 = 16'h0001; // 0x2526
	13'h1294: q1 = 16'h758e; // 0x2528
	13'h1295: q1 = 16'h670c; // 0x252a
	13'h1296: q1 = 16'h33c7; // 0x252c
	13'h1297: q1 = 16'h0001; // 0x252e
	13'h1298: q1 = 16'h7fa6; // 0x2530
	13'h1299: q1 = 16'h33c7; // 0x2532
	13'h129a: q1 = 16'h0001; // 0x2534
	13'h129b: q1 = 16'h8052; // 0x2536
	13'h129c: q1 = 16'h33fc; // 0x2538
	13'h129d: q1 = 16'h0001; // 0x253a
	13'h129e: q1 = 16'h0001; // 0x253c
	13'h129f: q1 = 16'h7f20; // 0x253e
	13'h12a0: q1 = 16'h3d7c; // 0x2540
	13'h12a1: q1 = 16'h002d; // 0x2542
	13'h12a2: q1 = 16'hfff2; // 0x2544
	13'h12a3: q1 = 16'h23fc; // 0x2546
	13'h12a4: q1 = 16'h0000; // 0x2548
	13'h12a5: q1 = 16'h003c; // 0x254a
	13'h12a6: q1 = 16'h0001; // 0x254c
	13'h12a7: q1 = 16'h7fac; // 0x254e
	13'h12a8: q1 = 16'h3d7c; // 0x2550
	13'h12a9: q1 = 16'h001e; // 0x2552
	13'h12aa: q1 = 16'hffe2; // 0x2554
	13'h12ab: q1 = 16'h2d79; // 0x2556
	13'h12ac: q1 = 16'h0000; // 0x2558
	13'h12ad: q1 = 16'hcca2; // 0x255a
	13'h12ae: q1 = 16'hffee; // 0x255c
	13'h12af: q1 = 16'h3d7c; // 0x255e
	13'h12b0: q1 = 16'h0001; // 0x2560
	13'h12b1: q1 = 16'hffe4; // 0x2562
	13'h12b2: q1 = 16'h3ebc; // 0x2564
	13'h12b3: q1 = 16'h0017; // 0x2566
	13'h12b4: q1 = 16'h4eb9; // 0x2568
	13'h12b5: q1 = 16'h0000; // 0x256a
	13'h12b6: q1 = 16'h8a22; // 0x256c
	13'h12b7: q1 = 16'h3ebc; // 0x256e
	13'h12b8: q1 = 16'h0018; // 0x2570
	13'h12b9: q1 = 16'h4eb9; // 0x2572
	13'h12ba: q1 = 16'h0000; // 0x2574
	13'h12bb: q1 = 16'h8a22; // 0x2576
	13'h12bc: q1 = 16'h4245; // 0x2578
	13'h12bd: q1 = 16'hba7c; // 0x257a
	13'h12be: q1 = 16'h001c; // 0x257c
	13'h12bf: q1 = 16'h6c3a; // 0x257e
	13'h12c0: q1 = 16'h3ebc; // 0x2580
	13'h12c1: q1 = 16'h003e; // 0x2582
	13'h12c2: q1 = 16'h3f05; // 0x2584
	13'h12c3: q1 = 16'h0657; // 0x2586
	13'h12c4: q1 = 16'h0041; // 0x2588
	13'h12c5: q1 = 16'h3005; // 0x258a
	13'h12c6: q1 = 16'h48c0; // 0x258c
	13'h12c7: q1 = 16'hd0bc; // 0x258e
	13'h12c8: q1 = 16'h0000; // 0x2590
	13'h12c9: q1 = 16'hcc86; // 0x2592
	13'h12ca: q1 = 16'h2040; // 0x2594
	13'h12cb: q1 = 16'h1010; // 0x2596
	13'h12cc: q1 = 16'h4880; // 0x2598
	13'h12cd: q1 = 16'h3f00; // 0x259a
	13'h12ce: q1 = 16'h3005; // 0x259c
	13'h12cf: q1 = 16'h48c0; // 0x259e
	13'h12d0: q1 = 16'hd0bc; // 0x25a0
	13'h12d1: q1 = 16'h0000; // 0x25a2
	13'h12d2: q1 = 16'hcc6a; // 0x25a4
	13'h12d3: q1 = 16'h2040; // 0x25a6
	13'h12d4: q1 = 16'h1010; // 0x25a8
	13'h12d5: q1 = 16'h4880; // 0x25aa
	13'h12d6: q1 = 16'h3f00; // 0x25ac
	13'h12d7: q1 = 16'h4eb9; // 0x25ae
	13'h12d8: q1 = 16'h0000; // 0x25b0
	13'h12d9: q1 = 16'h3d18; // 0x25b2
	13'h12da: q1 = 16'h5c4f; // 0x25b4
	13'h12db: q1 = 16'h5245; // 0x25b6
	13'h12dc: q1 = 16'h60c0; // 0x25b8
	13'h12dd: q1 = 16'h2eb9; // 0x25ba
	13'h12de: q1 = 16'h0000; // 0x25bc
	13'h12df: q1 = 16'hcca6; // 0x25be
	13'h12e0: q1 = 16'h4eb9; // 0x25c0
	13'h12e1: q1 = 16'h0000; // 0x25c2
	13'h12e2: q1 = 16'h3a7c; // 0x25c4
	13'h12e3: q1 = 16'h4eb9; // 0x25c6
	13'h12e4: q1 = 16'h0000; // 0x25c8
	13'h12e5: q1 = 16'h8680; // 0x25ca
	13'h12e6: q1 = 16'h4eb9; // 0x25cc
	13'h12e7: q1 = 16'h0000; // 0x25ce
	13'h12e8: q1 = 16'h47e8; // 0x25d0
	13'h12e9: q1 = 16'h200d; // 0x25d2
	13'h12ea: q1 = 16'h5080; // 0x25d4
	13'h12eb: q1 = 16'h2e80; // 0x25d6
	13'h12ec: q1 = 16'h200e; // 0x25d8
	13'h12ed: q1 = 16'hd0bc; // 0x25da
	13'h12ee: q1 = 16'hffff; // 0x25dc
	13'h12ef: q1 = 16'hffc0; // 0x25de
	13'h12f0: q1 = 16'h2f00; // 0x25e0
	13'h12f1: q1 = 16'h4eb9; // 0x25e2
	13'h12f2: q1 = 16'h0000; // 0x25e4
	13'h12f3: q1 = 16'h0750; // 0x25e6
	13'h12f4: q1 = 16'h4a9f; // 0x25e8
	13'h12f5: q1 = 16'h3ebc; // 0x25ea
	13'h12f6: q1 = 16'h003a; // 0x25ec
	13'h12f7: q1 = 16'h4267; // 0x25ee
	13'h12f8: q1 = 16'h3f3c; // 0x25f0
	13'h12f9: q1 = 16'hffeb; // 0x25f2
	13'h12fa: q1 = 16'h3f3c; // 0x25f4
	13'h12fb: q1 = 16'h0016; // 0x25f6
	13'h12fc: q1 = 16'h200e; // 0x25f8
	13'h12fd: q1 = 16'hd0bc; // 0x25fa
	13'h12fe: q1 = 16'hffff; // 0x25fc
	13'h12ff: q1 = 16'hffc0; // 0x25fe
	13'h1300: q1 = 16'h2f00; // 0x2600
	13'h1301: q1 = 16'h4eb9; // 0x2602
	13'h1302: q1 = 16'h0000; // 0x2604
	13'h1303: q1 = 16'h026c; // 0x2606
	13'h1304: q1 = 16'hdefc; // 0x2608
	13'h1305: q1 = 16'h000a; // 0x260a
	13'h1306: q1 = 16'h3ebc; // 0x260c
	13'h1307: q1 = 16'h0020; // 0x260e
	13'h1308: q1 = 16'h200e; // 0x2610
	13'h1309: q1 = 16'hd0bc; // 0x2612
	13'h130a: q1 = 16'hffff; // 0x2614
	13'h130b: q1 = 16'hfff4; // 0x2616
	13'h130c: q1 = 16'h2f00; // 0x2618
	13'h130d: q1 = 16'h200e; // 0x261a
	13'h130e: q1 = 16'hd0bc; // 0x261c
	13'h130f: q1 = 16'hffff; // 0x261e
	13'h1310: q1 = 16'hffec; // 0x2620
	13'h1311: q1 = 16'h2f00; // 0x2622
	13'h1312: q1 = 16'h3f15; // 0x2624
	13'h1313: q1 = 16'h4eb9; // 0x2626
	13'h1314: q1 = 16'h0000; // 0x2628
	13'h1315: q1 = 16'h1402; // 0x262a
	13'h1316: q1 = 16'hdefc; // 0x262c
	13'h1317: q1 = 16'h000a; // 0x262e
	13'h1318: q1 = 16'h0c6e; // 0x2630
	13'h1319: q1 = 16'h0001; // 0x2632
	13'h131a: q1 = 16'hffec; // 0x2634
	13'h131b: q1 = 16'h6608; // 0x2636
	13'h131c: q1 = 16'h3d7c; // 0x2638
	13'h131d: q1 = 16'h00e9; // 0x263a
	13'h131e: q1 = 16'hffea; // 0x263c
	13'h131f: q1 = 16'h6016; // 0x263e
	13'h1320: q1 = 16'h0c6e; // 0x2640
	13'h1321: q1 = 16'h0002; // 0x2642
	13'h1322: q1 = 16'hffec; // 0x2644
	13'h1323: q1 = 16'h6608; // 0x2646
	13'h1324: q1 = 16'h3d7c; // 0x2648
	13'h1325: q1 = 16'h00e1; // 0x264a
	13'h1326: q1 = 16'hffea; // 0x264c
	13'h1327: q1 = 16'h6006; // 0x264e
	13'h1328: q1 = 16'h3d7c; // 0x2650
	13'h1329: q1 = 16'h00d9; // 0x2652
	13'h132a: q1 = 16'hffea; // 0x2654
	13'h132b: q1 = 16'h3ebc; // 0x2656
	13'h132c: q1 = 16'h0020; // 0x2658
	13'h132d: q1 = 16'h3f2e; // 0x265a
	13'h132e: q1 = 16'hffea; // 0x265c
	13'h132f: q1 = 16'h3f3c; // 0x265e
	13'h1330: q1 = 16'h0016; // 0x2660
	13'h1331: q1 = 16'h3f3c; // 0x2662
	13'h1332: q1 = 16'h0017; // 0x2664
	13'h1333: q1 = 16'h4eb9; // 0x2666
	13'h1334: q1 = 16'h0000; // 0x2668
	13'h1335: q1 = 16'h3d18; // 0x266a
	13'h1336: q1 = 16'h5c4f; // 0x266c
	13'h1337: q1 = 16'h3ebc; // 0x266e
	13'h1338: q1 = 16'h0021; // 0x2670
	13'h1339: q1 = 16'h3f39; // 0x2672
	13'h133a: q1 = 16'h0000; // 0x2674
	13'h133b: q1 = 16'hca9c; // 0x2676
	13'h133c: q1 = 16'h3f3c; // 0x2678
	13'h133d: q1 = 16'h0015; // 0x267a
	13'h133e: q1 = 16'h3f3c; // 0x267c
	13'h133f: q1 = 16'h0017; // 0x267e
	13'h1340: q1 = 16'h4eb9; // 0x2680
	13'h1341: q1 = 16'h0000; // 0x2682
	13'h1342: q1 = 16'h3d18; // 0x2684
	13'h1343: q1 = 16'h5c4f; // 0x2686
	13'h1344: q1 = 16'h4245; // 0x2688
	13'h1345: q1 = 16'h3d7c; // 0x268a
	13'h1346: q1 = 16'h005c; // 0x268c
	13'h1347: q1 = 16'hfffc; // 0x268e
	13'h1348: q1 = 16'h3d7c; // 0x2690
	13'h1349: q1 = 16'h005c; // 0x2692
	13'h134a: q1 = 16'hffea; // 0x2694
	13'h134b: q1 = 16'h3d7c; // 0x2696
	13'h134c: q1 = 16'h0020; // 0x2698
	13'h134d: q1 = 16'hfffa; // 0x269a
	13'h134e: q1 = 16'h426e; // 0x269c
	13'h134f: q1 = 16'hffbe; // 0x269e
	13'h1350: q1 = 16'h7c08; // 0x26a0
	13'h1351: q1 = 16'hbc7c; // 0x26a2
	13'h1352: q1 = 16'h000a; // 0x26a4
	13'h1353: q1 = 16'h6e1a; // 0x26a6
	13'h1354: q1 = 16'h3ebc; // 0x26a8
	13'h1355: q1 = 16'h003c; // 0x26aa
	13'h1356: q1 = 16'h3f3c; // 0x26ac
	13'h1357: q1 = 16'h005c; // 0x26ae
	13'h1358: q1 = 16'h3f3c; // 0x26b0
	13'h1359: q1 = 16'h0016; // 0x26b2
	13'h135a: q1 = 16'h3f06; // 0x26b4
	13'h135b: q1 = 16'h4eb9; // 0x26b6
	13'h135c: q1 = 16'h0000; // 0x26b8
	13'h135d: q1 = 16'h3d18; // 0x26ba
	13'h135e: q1 = 16'h5c4f; // 0x26bc
	13'h135f: q1 = 16'h5246; // 0x26be
	13'h1360: q1 = 16'h60e0; // 0x26c0
	13'h1361: q1 = 16'h3d7c; // 0x26c2
	13'h1362: q1 = 16'h001b; // 0x26c4
	13'h1363: q1 = 16'hfffe; // 0x26c6
	13'h1364: q1 = 16'h23fc; // 0x26c8
	13'h1365: q1 = 16'h0000; // 0x26ca
	13'h1366: q1 = 16'h0002; // 0x26cc
	13'h1367: q1 = 16'h0001; // 0x26ce
	13'h1368: q1 = 16'h7fc2; // 0x26d0
	13'h1369: q1 = 16'h4ab9; // 0x26d2
	13'h136a: q1 = 16'h0001; // 0x26d4
	13'h136b: q1 = 16'h7fac; // 0x26d6
	13'h136c: q1 = 16'h660e; // 0x26d8
	13'h136d: q1 = 16'h536e; // 0x26da
	13'h136e: q1 = 16'hffe2; // 0x26dc
	13'h136f: q1 = 16'h23fc; // 0x26de
	13'h1370: q1 = 16'h0000; // 0x26e0
	13'h1371: q1 = 16'h003c; // 0x26e2
	13'h1372: q1 = 16'h0001; // 0x26e4
	13'h1373: q1 = 16'h7fac; // 0x26e6
	13'h1374: q1 = 16'h3ebc; // 0x26e8
	13'h1375: q1 = 16'h000e; // 0x26ea
	13'h1376: q1 = 16'h200e; // 0x26ec
	13'h1377: q1 = 16'hd0bc; // 0x26ee
	13'h1378: q1 = 16'hffff; // 0x26f0
	13'h1379: q1 = 16'hffc0; // 0x26f2
	13'h137a: q1 = 16'h2f00; // 0x26f4
	13'h137b: q1 = 16'h4eb9; // 0x26f6
	13'h137c: q1 = 16'h0000; // 0x26f8
	13'h137d: q1 = 16'h78f6; // 0x26fa
	13'h137e: q1 = 16'h4a9f; // 0x26fc
	13'h137f: q1 = 16'h0c6e; // 0x26fe
	13'h1380: q1 = 16'h000a; // 0x2700
	13'h1381: q1 = 16'hffe2; // 0x2702
	13'h1382: q1 = 16'h6c18; // 0x2704
	13'h1383: q1 = 16'h2ebc; // 0x2706
	13'h1384: q1 = 16'h0000; // 0x2708
	13'h1385: q1 = 16'hccaa; // 0x270a
	13'h1386: q1 = 16'h200e; // 0x270c
	13'h1387: q1 = 16'hd0bc; // 0x270e
	13'h1388: q1 = 16'hffff; // 0x2710
	13'h1389: q1 = 16'hffc0; // 0x2712
	13'h138a: q1 = 16'h2f00; // 0x2714
	13'h138b: q1 = 16'h4eb9; // 0x2716
	13'h138c: q1 = 16'h0000; // 0x2718
	13'h138d: q1 = 16'h0770; // 0x271a
	13'h138e: q1 = 16'h4a9f; // 0x271c
	13'h138f: q1 = 16'h200e; // 0x271e
	13'h1390: q1 = 16'hd0bc; // 0x2720
	13'h1391: q1 = 16'hffff; // 0x2722
	13'h1392: q1 = 16'hffc0; // 0x2724
	13'h1393: q1 = 16'h2e80; // 0x2726
	13'h1394: q1 = 16'h3f2e; // 0x2728
	13'h1395: q1 = 16'hffe2; // 0x272a
	13'h1396: q1 = 16'h4eb9; // 0x272c
	13'h1397: q1 = 16'h0000; // 0x272e
	13'h1398: q1 = 16'h0798; // 0x2730
	13'h1399: q1 = 16'h4a5f; // 0x2732
	13'h139a: q1 = 16'h3ebc; // 0x2734
	13'h139b: q1 = 16'h0031; // 0x2736
	13'h139c: q1 = 16'h4267; // 0x2738
	13'h139d: q1 = 16'h3f3c; // 0x273a
	13'h139e: q1 = 16'h0064; // 0x273c
	13'h139f: q1 = 16'h3f3c; // 0x273e
	13'h13a0: q1 = 16'h000c; // 0x2740
	13'h13a1: q1 = 16'h200e; // 0x2742
	13'h13a2: q1 = 16'hd0bc; // 0x2744
	13'h13a3: q1 = 16'hffff; // 0x2746
	13'h13a4: q1 = 16'hffc0; // 0x2748
	13'h13a5: q1 = 16'h2f00; // 0x274a
	13'h13a6: q1 = 16'h4eb9; // 0x274c
	13'h13a7: q1 = 16'h0000; // 0x274e
	13'h13a8: q1 = 16'h026c; // 0x2750
	13'h13a9: q1 = 16'hdefc; // 0x2752
	13'h13aa: q1 = 16'h000a; // 0x2754
	13'h13ab: q1 = 16'h4a6e; // 0x2756
	13'h13ac: q1 = 16'hffe2; // 0x2758
	13'h13ad: q1 = 16'h6700; // 0x275a
	13'h13ae: q1 = 16'h035e; // 0x275c
	13'h13af: q1 = 16'h4a79; // 0x275e
	13'h13b0: q1 = 16'h0001; // 0x2760
	13'h13b1: q1 = 16'h7f5e; // 0x2762
	13'h13b2: q1 = 16'h6600; // 0x2764
	13'h13b3: q1 = 16'h0354; // 0x2766
	13'h13b4: q1 = 16'h3ebc; // 0x2768
	13'h13b5: q1 = 16'h0033; // 0x276a
	13'h13b6: q1 = 16'h200e; // 0x276c
	13'h13b7: q1 = 16'hd0bc; // 0x276e
	13'h13b8: q1 = 16'hffff; // 0x2770
	13'h13b9: q1 = 16'hffc0; // 0x2772
	13'h13ba: q1 = 16'h2f00; // 0x2774
	13'h13bb: q1 = 16'h4eb9; // 0x2776
	13'h13bc: q1 = 16'h0000; // 0x2778
	13'h13bd: q1 = 16'h78f6; // 0x277a
	13'h13be: q1 = 16'h4a9f; // 0x277c
	13'h13bf: q1 = 16'h200e; // 0x277e
	13'h13c0: q1 = 16'hd0bc; // 0x2780
	13'h13c1: q1 = 16'hffff; // 0x2782
	13'h13c2: q1 = 16'hffc0; // 0x2784
	13'h13c3: q1 = 16'h2e80; // 0x2786
	13'h13c4: q1 = 16'h3f07; // 0x2788
	13'h13c5: q1 = 16'h5257; // 0x278a
	13'h13c6: q1 = 16'h4eb9; // 0x278c
	13'h13c7: q1 = 16'h0000; // 0x278e
	13'h13c8: q1 = 16'h0798; // 0x2790
	13'h13c9: q1 = 16'h4a5f; // 0x2792
	13'h13ca: q1 = 16'h0c79; // 0x2794
	13'h13cb: q1 = 16'h0002; // 0x2796
	13'h13cc: q1 = 16'h0001; // 0x2798
	13'h13cd: q1 = 16'h758c; // 0x279a
	13'h13ce: q1 = 16'h6718; // 0x279c
	13'h13cf: q1 = 16'h2ebc; // 0x279e
	13'h13d0: q1 = 16'h0000; // 0x27a0
	13'h13d1: q1 = 16'hccac; // 0x27a2
	13'h13d2: q1 = 16'h200e; // 0x27a4
	13'h13d3: q1 = 16'hd0bc; // 0x27a6
	13'h13d4: q1 = 16'hffff; // 0x27a8
	13'h13d5: q1 = 16'hffc0; // 0x27aa
	13'h13d6: q1 = 16'h2f00; // 0x27ac
	13'h13d7: q1 = 16'h4eb9; // 0x27ae
	13'h13d8: q1 = 16'h0000; // 0x27b0
	13'h13d9: q1 = 16'h0770; // 0x27b2
	13'h13da: q1 = 16'h4a9f; // 0x27b4
	13'h13db: q1 = 16'h2ebc; // 0x27b6
	13'h13dc: q1 = 16'h0000; // 0x27b8
	13'h13dd: q1 = 16'hccae; // 0x27ba
	13'h13de: q1 = 16'h200e; // 0x27bc
	13'h13df: q1 = 16'hd0bc; // 0x27be
	13'h13e0: q1 = 16'hffff; // 0x27c0
	13'h13e1: q1 = 16'hffc0; // 0x27c2
	13'h13e2: q1 = 16'h2f00; // 0x27c4
	13'h13e3: q1 = 16'h4eb9; // 0x27c6
	13'h13e4: q1 = 16'h0000; // 0x27c8
	13'h13e5: q1 = 16'h0770; // 0x27ca
	13'h13e6: q1 = 16'h4a9f; // 0x27cc
	13'h13e7: q1 = 16'h3eae; // 0x27ce
	13'h13e8: q1 = 16'hfff2; // 0x27d0
	13'h13e9: q1 = 16'h4267; // 0x27d2
	13'h13ea: q1 = 16'h3f3c; // 0x27d4
	13'h13eb: q1 = 16'h0064; // 0x27d6
	13'h13ec: q1 = 16'h3f3c; // 0x27d8
	13'h13ed: q1 = 16'h001f; // 0x27da
	13'h13ee: q1 = 16'h200e; // 0x27dc
	13'h13ef: q1 = 16'hd0bc; // 0x27de
	13'h13f0: q1 = 16'hffff; // 0x27e0
	13'h13f1: q1 = 16'hffc0; // 0x27e2
	13'h13f2: q1 = 16'h2f00; // 0x27e4
	13'h13f3: q1 = 16'h4eb9; // 0x27e6
	13'h13f4: q1 = 16'h0000; // 0x27e8
	13'h13f5: q1 = 16'h026c; // 0x27ea
	13'h13f6: q1 = 16'hdefc; // 0x27ec
	13'h13f7: q1 = 16'h000a; // 0x27ee
	13'h13f8: q1 = 16'h526e; // 0x27f0
	13'h13f9: q1 = 16'hfff2; // 0x27f2
	13'h13fa: q1 = 16'h0c6e; // 0x27f4
	13'h13fb: q1 = 16'h003f; // 0x27f6
	13'h13fc: q1 = 16'hfff2; // 0x27f8
	13'h13fd: q1 = 16'h6f06; // 0x27fa
	13'h13fe: q1 = 16'h3d7c; // 0x27fc
	13'h13ff: q1 = 16'h002d; // 0x27fe
	13'h1400: q1 = 16'hfff2; // 0x2800
	13'h1401: q1 = 16'h4a79; // 0x2802
	13'h1402: q1 = 16'h0001; // 0x2804
	13'h1403: q1 = 16'h7fca; // 0x2806
	13'h1404: q1 = 16'h6700; // 0x2808
	13'h1405: q1 = 16'h00ac; // 0x280a
	13'h1406: q1 = 16'h4a6e; // 0x280c
	13'h1407: q1 = 16'hffe4; // 0x280e
	13'h1408: q1 = 16'h6600; // 0x2810
	13'h1409: q1 = 16'h00a4; // 0x2812
	13'h140a: q1 = 16'h3d7c; // 0x2814
	13'h140b: q1 = 16'h0001; // 0x2816
	13'h140c: q1 = 16'hffe4; // 0x2818
	13'h140d: q1 = 16'h0c6e; // 0x281a
	13'h140e: q1 = 16'h001a; // 0x281c
	13'h140f: q1 = 16'hfffe; // 0x281e
	13'h1410: q1 = 16'h6608; // 0x2820
	13'h1411: q1 = 16'h3d7c; // 0x2822
	13'h1412: q1 = 16'h003c; // 0x2824
	13'h1413: q1 = 16'hffe8; // 0x2826
	13'h1414: q1 = 16'h6006; // 0x2828
	13'h1415: q1 = 16'h3d7c; // 0x282a
	13'h1416: q1 = 16'h003a; // 0x282c
	13'h1417: q1 = 16'hffe8; // 0x282e
	13'h1418: q1 = 16'h3eae; // 0x2830
	13'h1419: q1 = 16'hffe8; // 0x2832
	13'h141a: q1 = 16'h3f2e; // 0x2834
	13'h141b: q1 = 16'hffea; // 0x2836
	13'h141c: q1 = 16'h3f3c; // 0x2838
	13'h141d: q1 = 16'h0016; // 0x283a
	13'h141e: q1 = 16'h3f05; // 0x283c
	13'h141f: q1 = 16'h5057; // 0x283e
	13'h1420: q1 = 16'h4eb9; // 0x2840
	13'h1421: q1 = 16'h0000; // 0x2842
	13'h1422: q1 = 16'h3d18; // 0x2844
	13'h1423: q1 = 16'h5c4f; // 0x2846
	13'h1424: q1 = 16'h0c6e; // 0x2848
	13'h1425: q1 = 16'h001a; // 0x284a
	13'h1426: q1 = 16'hfffe; // 0x284c
	13'h1427: q1 = 16'h664a; // 0x284e
	13'h1428: q1 = 16'h4a45; // 0x2850
	13'h1429: q1 = 16'h6f40; // 0x2852
	13'h142a: q1 = 16'h5345; // 0x2854
	13'h142b: q1 = 16'h200e; // 0x2856
	13'h142c: q1 = 16'hd0bc; // 0x2858
	13'h142d: q1 = 16'hffff; // 0x285a
	13'h142e: q1 = 16'hffe8; // 0x285c
	13'h142f: q1 = 16'h2e80; // 0x285e
	13'h1430: q1 = 16'h200e; // 0x2860
	13'h1431: q1 = 16'hd0bc; // 0x2862
	13'h1432: q1 = 16'hffff; // 0x2864
	13'h1433: q1 = 16'hffe6; // 0x2866
	13'h1434: q1 = 16'h2f00; // 0x2868
	13'h1435: q1 = 16'h3f3c; // 0x286a
	13'h1436: q1 = 16'h0016; // 0x286c
	13'h1437: q1 = 16'h3f05; // 0x286e
	13'h1438: q1 = 16'h5057; // 0x2870
	13'h1439: q1 = 16'h4eb9; // 0x2872
	13'h143a: q1 = 16'h0000; // 0x2874
	13'h143b: q1 = 16'h3dbe; // 0x2876
	13'h143c: q1 = 16'hbf8f; // 0x2878
	13'h143d: q1 = 16'h3ebc; // 0x287a
	13'h143e: q1 = 16'h003c; // 0x287c
	13'h143f: q1 = 16'h3f2e; // 0x287e
	13'h1440: q1 = 16'hffe6; // 0x2880
	13'h1441: q1 = 16'h3f3c; // 0x2882
	13'h1442: q1 = 16'h0016; // 0x2884
	13'h1443: q1 = 16'h3f05; // 0x2886
	13'h1444: q1 = 16'h5057; // 0x2888
	13'h1445: q1 = 16'h4eb9; // 0x288a
	13'h1446: q1 = 16'h0000; // 0x288c
	13'h1447: q1 = 16'h3d18; // 0x288e
	13'h1448: q1 = 16'h5c4f; // 0x2890
	13'h1449: q1 = 16'h6004; // 0x2892
	13'h144a: q1 = 16'h526e; // 0x2894
	13'h144b: q1 = 16'hffbe; // 0x2896
	13'h144c: q1 = 16'h6012; // 0x2898
	13'h144d: q1 = 16'h3005; // 0x289a
	13'h144e: q1 = 16'he340; // 0x289c
	13'h144f: q1 = 16'h48c0; // 0x289e
	13'h1450: q1 = 16'hd08e; // 0x28a0
	13'h1451: q1 = 16'h2040; // 0x28a2
	13'h1452: q1 = 16'h316e; // 0x28a4
	13'h1453: q1 = 16'hfffa; // 0x28a6
	13'h1454: q1 = 16'hfff4; // 0x28a8
	13'h1455: q1 = 16'h5245; // 0x28aa
	13'h1456: q1 = 16'hba7c; // 0x28ac
	13'h1457: q1 = 16'h0003; // 0x28ae
	13'h1458: q1 = 16'h6700; // 0x28b0
	13'h1459: q1 = 16'h0194; // 0x28b2
	13'h145a: q1 = 16'h6012; // 0x28b4
	13'h145b: q1 = 16'h4a6e; // 0x28b6
	13'h145c: q1 = 16'hffe4; // 0x28b8
	13'h145d: q1 = 16'h670c; // 0x28ba
	13'h145e: q1 = 16'h4a79; // 0x28bc
	13'h145f: q1 = 16'h0001; // 0x28be
	13'h1460: q1 = 16'h7fca; // 0x28c0
	13'h1461: q1 = 16'h6604; // 0x28c2
	13'h1462: q1 = 16'h426e; // 0x28c4
	13'h1463: q1 = 16'hffe4; // 0x28c6
	13'h1464: q1 = 16'h4eb9; // 0x28c8
	13'h1465: q1 = 16'h0000; // 0x28ca
	13'h1466: q1 = 16'h4820; // 0x28cc
	13'h1467: q1 = 16'h4eb9; // 0x28ce
	13'h1468: q1 = 16'h0000; // 0x28d0
	13'h1469: q1 = 16'h3434; // 0x28d2
	13'h146a: q1 = 16'h4246; // 0x28d4
	13'h146b: q1 = 16'hbc7c; // 0x28d6
	13'h146c: q1 = 16'h001c; // 0x28d8
	13'h146d: q1 = 16'h6c00; // 0x28da
	13'h146e: q1 = 16'h014a; // 0x28dc
	13'h146f: q1 = 16'h3006; // 0x28de
	13'h1470: q1 = 16'h48c0; // 0x28e0
	13'h1471: q1 = 16'hd0bc; // 0x28e2
	13'h1472: q1 = 16'h0000; // 0x28e4
	13'h1473: q1 = 16'hcc6a; // 0x28e6
	13'h1474: q1 = 16'h2040; // 0x28e8
	13'h1475: q1 = 16'h1810; // 0x28ea
	13'h1476: q1 = 16'h4884; // 0x28ec
	13'h1477: q1 = 16'h4280; // 0x28ee
	13'h1478: q1 = 16'h700a; // 0x28f0
	13'h1479: q1 = 16'he164; // 0x28f2
	13'h147a: q1 = 16'h3006; // 0x28f4
	13'h147b: q1 = 16'h48c0; // 0x28f6
	13'h147c: q1 = 16'hd0bc; // 0x28f8
	13'h147d: q1 = 16'h0000; // 0x28fa
	13'h147e: q1 = 16'hcc86; // 0x28fc
	13'h147f: q1 = 16'h2040; // 0x28fe
	13'h1480: q1 = 16'h1610; // 0x2900
	13'h1481: q1 = 16'h4883; // 0x2902
	13'h1482: q1 = 16'h4280; // 0x2904
	13'h1483: q1 = 16'h700a; // 0x2906
	13'h1484: q1 = 16'he163; // 0x2908
	13'h1485: q1 = 16'h200e; // 0x290a
	13'h1486: q1 = 16'hd0bc; // 0x290c
	13'h1487: q1 = 16'hffff; // 0x290e
	13'h1488: q1 = 16'hffec; // 0x2910
	13'h1489: q1 = 16'h2e80; // 0x2912
	13'h148a: q1 = 16'h200e; // 0x2914
	13'h148b: q1 = 16'hd0bc; // 0x2916
	13'h148c: q1 = 16'hffff; // 0x2918
	13'h148d: q1 = 16'hffec; // 0x291a
	13'h148e: q1 = 16'h2f00; // 0x291c
	13'h148f: q1 = 16'h200e; // 0x291e
	13'h1490: q1 = 16'hd0bc; // 0x2920
	13'h1491: q1 = 16'hffff; // 0x2922
	13'h1492: q1 = 16'hffec; // 0x2924
	13'h1493: q1 = 16'h2f00; // 0x2926
	13'h1494: q1 = 16'h200e; // 0x2928
	13'h1495: q1 = 16'hd0bc; // 0x292a
	13'h1496: q1 = 16'hffff; // 0x292c
	13'h1497: q1 = 16'hffec; // 0x292e
	13'h1498: q1 = 16'h2f00; // 0x2930
	13'h1499: q1 = 16'h2f2e; // 0x2932
	13'h149a: q1 = 16'hffee; // 0x2934
	13'h149b: q1 = 16'h3f03; // 0x2936
	13'h149c: q1 = 16'h0657; // 0x2938
	13'h149d: q1 = 16'hfe00; // 0x293a
	13'h149e: q1 = 16'h3f04; // 0x293c
	13'h149f: q1 = 16'h0657; // 0x293e
	13'h14a0: q1 = 16'hfe00; // 0x2940
	13'h14a1: q1 = 16'h4eb9; // 0x2942
	13'h14a2: q1 = 16'h0000; // 0x2944
	13'h14a3: q1 = 16'h36d8; // 0x2946
	13'h14a4: q1 = 16'hdefc; // 0x2948
	13'h14a5: q1 = 16'h0014; // 0x294a
	13'h14a6: q1 = 16'h4a80; // 0x294c
	13'h14a7: q1 = 16'h6700; // 0x294e
	13'h14a8: q1 = 16'h00d0; // 0x2950
	13'h14a9: q1 = 16'h302e; // 0x2952
	13'h14aa: q1 = 16'hfffe; // 0x2954
	13'h14ab: q1 = 16'hb046; // 0x2956
	13'h14ac: q1 = 16'h677c; // 0x2958
	13'h14ad: q1 = 16'h3ebc; // 0x295a
	13'h14ae: q1 = 16'h003e; // 0x295c
	13'h14af: q1 = 16'h3f2e; // 0x295e
	13'h14b0: q1 = 16'hfffc; // 0x2960
	13'h14b1: q1 = 16'h302e; // 0x2962
	13'h14b2: q1 = 16'hfffe; // 0x2964
	13'h14b3: q1 = 16'h48c0; // 0x2966
	13'h14b4: q1 = 16'hd0bc; // 0x2968
	13'h14b5: q1 = 16'h0000; // 0x296a
	13'h14b6: q1 = 16'hcc86; // 0x296c
	13'h14b7: q1 = 16'h2040; // 0x296e
	13'h14b8: q1 = 16'h1010; // 0x2970
	13'h14b9: q1 = 16'h4880; // 0x2972
	13'h14ba: q1 = 16'h3f00; // 0x2974
	13'h14bb: q1 = 16'h302e; // 0x2976
	13'h14bc: q1 = 16'hfffe; // 0x2978
	13'h14bd: q1 = 16'h48c0; // 0x297a
	13'h14be: q1 = 16'hd0bc; // 0x297c
	13'h14bf: q1 = 16'h0000; // 0x297e
	13'h14c0: q1 = 16'hcc6a; // 0x2980
	13'h14c1: q1 = 16'h2040; // 0x2982
	13'h14c2: q1 = 16'h1010; // 0x2984
	13'h14c3: q1 = 16'h4880; // 0x2986
	13'h14c4: q1 = 16'h3f00; // 0x2988
	13'h14c5: q1 = 16'h4eb9; // 0x298a
	13'h14c6: q1 = 16'h0000; // 0x298c
	13'h14c7: q1 = 16'h3d18; // 0x298e
	13'h14c8: q1 = 16'h5c4f; // 0x2990
	13'h14c9: q1 = 16'h200e; // 0x2992
	13'h14ca: q1 = 16'hd0bc; // 0x2994
	13'h14cb: q1 = 16'hffff; // 0x2996
	13'h14cc: q1 = 16'hffe8; // 0x2998
	13'h14cd: q1 = 16'h2e80; // 0x299a
	13'h14ce: q1 = 16'h200e; // 0x299c
	13'h14cf: q1 = 16'hd0bc; // 0x299e
	13'h14d0: q1 = 16'hffff; // 0x29a0
	13'h14d1: q1 = 16'hfffc; // 0x29a2
	13'h14d2: q1 = 16'h2f00; // 0x29a4
	13'h14d3: q1 = 16'h3f03; // 0x29a6
	13'h14d4: q1 = 16'h3f04; // 0x29a8
	13'h14d5: q1 = 16'h4eb9; // 0x29aa
	13'h14d6: q1 = 16'h0000; // 0x29ac
	13'h14d7: q1 = 16'h3dbe; // 0x29ae
	13'h14d8: q1 = 16'hbf8f; // 0x29b0
	13'h14d9: q1 = 16'h3ebc; // 0x29b2
	13'h14da: q1 = 16'h003c; // 0x29b4
	13'h14db: q1 = 16'h3f2e; // 0x29b6
	13'h14dc: q1 = 16'hfffc; // 0x29b8
	13'h14dd: q1 = 16'h3003; // 0x29ba
	13'h14de: q1 = 16'h4281; // 0x29bc
	13'h14df: q1 = 16'h720a; // 0x29be
	13'h14e0: q1 = 16'he260; // 0x29c0
	13'h14e1: q1 = 16'h3f00; // 0x29c2
	13'h14e2: q1 = 16'h3004; // 0x29c4
	13'h14e3: q1 = 16'h4281; // 0x29c6
	13'h14e4: q1 = 16'h720a; // 0x29c8
	13'h14e5: q1 = 16'he260; // 0x29ca
	13'h14e6: q1 = 16'h3f00; // 0x29cc
	13'h14e7: q1 = 16'h4eb9; // 0x29ce
	13'h14e8: q1 = 16'h0000; // 0x29d0
	13'h14e9: q1 = 16'h3d18; // 0x29d2
	13'h14ea: q1 = 16'h5c4f; // 0x29d4
	13'h14eb: q1 = 16'h3d6e; // 0x29d6
	13'h14ec: q1 = 16'hfffc; // 0x29d8
	13'h14ed: q1 = 16'hffea; // 0x29da
	13'h14ee: q1 = 16'hbc7c; // 0x29dc
	13'h14ef: q1 = 16'h001a; // 0x29de
	13'h14f0: q1 = 16'h6606; // 0x29e0
	13'h14f1: q1 = 16'h3d7c; // 0x29e2
	13'h14f2: q1 = 16'h005c; // 0x29e4
	13'h14f3: q1 = 16'hffea; // 0x29e6
	13'h14f4: q1 = 16'h4a6e; // 0x29e8
	13'h14f5: q1 = 16'hffe4; // 0x29ea
	13'h14f6: q1 = 16'h6618; // 0x29ec
	13'h14f7: q1 = 16'h3ebc; // 0x29ee
	13'h14f8: q1 = 16'h003c; // 0x29f0
	13'h14f9: q1 = 16'h3f2e; // 0x29f2
	13'h14fa: q1 = 16'hffea; // 0x29f4
	13'h14fb: q1 = 16'h3f3c; // 0x29f6
	13'h14fc: q1 = 16'h0016; // 0x29f8
	13'h14fd: q1 = 16'h3f05; // 0x29fa
	13'h14fe: q1 = 16'h5057; // 0x29fc
	13'h14ff: q1 = 16'h4eb9; // 0x29fe
	13'h1500: q1 = 16'h0000; // 0x2a00
	13'h1501: q1 = 16'h3d18; // 0x2a02
	13'h1502: q1 = 16'h5c4f; // 0x2a04
	13'h1503: q1 = 16'h3d46; // 0x2a06
	13'h1504: q1 = 16'hfffe; // 0x2a08
	13'h1505: q1 = 16'h3d6e; // 0x2a0a
	13'h1506: q1 = 16'hfffc; // 0x2a0c
	13'h1507: q1 = 16'hfffa; // 0x2a0e
	13'h1508: q1 = 16'h0c6e; // 0x2a10
	13'h1509: q1 = 16'h005c; // 0x2a12
	13'h150a: q1 = 16'hfffa; // 0x2a14
	13'h150b: q1 = 16'h6606; // 0x2a16
	13'h150c: q1 = 16'h3d7c; // 0x2a18
	13'h150d: q1 = 16'h0020; // 0x2a1a
	13'h150e: q1 = 16'hfffa; // 0x2a1c
	13'h150f: q1 = 16'h6006; // 0x2a1e
	13'h1510: q1 = 16'h5246; // 0x2a20
	13'h1511: q1 = 16'h6000; // 0x2a22
	13'h1512: q1 = 16'hfeb2; // 0x2a24
	13'h1513: q1 = 16'h4ab9; // 0x2a26
	13'h1514: q1 = 16'h0001; // 0x2a28
	13'h1515: q1 = 16'h7fc2; // 0x2a2a
	13'h1516: q1 = 16'h6714; // 0x2a2c
	13'h1517: q1 = 16'h4a6e; // 0x2a2e
	13'h1518: q1 = 16'hffe2; // 0x2a30
	13'h1519: q1 = 16'h6700; // 0x2a32
	13'h151a: q1 = 16'h0086; // 0x2a34
	13'h151b: q1 = 16'h4a79; // 0x2a36
	13'h151c: q1 = 16'h0001; // 0x2a38
	13'h151d: q1 = 16'h7f5e; // 0x2a3a
	13'h151e: q1 = 16'h6600; // 0x2a3c
	13'h151f: q1 = 16'h007c; // 0x2a3e
	13'h1520: q1 = 16'h60e4; // 0x2a40
	13'h1521: q1 = 16'h6000; // 0x2a42
	13'h1522: q1 = 16'hfc84; // 0x2a44
	13'h1523: q1 = 16'h3c2d; // 0x2a46
	13'h1524: q1 = 16'h001e; // 0x2a48
	13'h1525: q1 = 16'h5346; // 0x2a4a
	13'h1526: q1 = 16'h0c6e; // 0x2a4c
	13'h1527: q1 = 16'h0007; // 0x2a4e
	13'h1528: q1 = 16'hffbe; // 0x2a50
	13'h1529: q1 = 16'h6638; // 0x2a52
	13'h152a: q1 = 16'h0c6e; // 0x2a54
	13'h152b: q1 = 16'h004a; // 0x2a56
	13'h152c: q1 = 16'hfff4; // 0x2a58
	13'h152d: q1 = 16'h6630; // 0x2a5a
	13'h152e: q1 = 16'h0c6e; // 0x2a5c
	13'h152f: q1 = 16'h0041; // 0x2a5e
	13'h1530: q1 = 16'hfff6; // 0x2a60
	13'h1531: q1 = 16'h6628; // 0x2a62
	13'h1532: q1 = 16'h0c6e; // 0x2a64
	13'h1533: q1 = 16'h0048; // 0x2a66
	13'h1534: q1 = 16'hfff8; // 0x2a68
	13'h1535: q1 = 16'h6620; // 0x2a6a
	13'h1536: q1 = 16'h4245; // 0x2a6c
	13'h1537: q1 = 16'hba7c; // 0x2a6e
	13'h1538: q1 = 16'h0003; // 0x2a70
	13'h1539: q1 = 16'h6c18; // 0x2a72
	13'h153a: q1 = 16'h3005; // 0x2a74
	13'h153b: q1 = 16'he340; // 0x2a76
	13'h153c: q1 = 16'h48c0; // 0x2a78
	13'h153d: q1 = 16'hd08e; // 0x2a7a
	13'h153e: q1 = 16'h2040; // 0x2a7c
	13'h153f: q1 = 16'h3205; // 0x2a7e
	13'h1540: q1 = 16'hd27c; // 0x2a80
	13'h1541: q1 = 16'h0072; // 0x2a82
	13'h1542: q1 = 16'h3141; // 0x2a84
	13'h1543: q1 = 16'hfff4; // 0x2a86
	13'h1544: q1 = 16'h5245; // 0x2a88
	13'h1545: q1 = 16'h60e2; // 0x2a8a
	13'h1546: q1 = 16'h4245; // 0x2a8c
	13'h1547: q1 = 16'hba7c; // 0x2a8e
	13'h1548: q1 = 16'h0003; // 0x2a90
	13'h1549: q1 = 16'h6c26; // 0x2a92
	13'h154a: q1 = 16'h3006; // 0x2a94
	13'h154b: q1 = 16'hc1fc; // 0x2a96
	13'h154c: q1 = 16'h0003; // 0x2a98
	13'h154d: q1 = 16'hd045; // 0x2a9a
	13'h154e: q1 = 16'h48c0; // 0x2a9c
	13'h154f: q1 = 16'hd0bc; // 0x2a9e
	13'h1550: q1 = 16'h0001; // 0x2aa0
	13'h1551: q1 = 16'h7ba8; // 0x2aa2
	13'h1552: q1 = 16'h2040; // 0x2aa4
	13'h1553: q1 = 16'h3205; // 0x2aa6
	13'h1554: q1 = 16'he341; // 0x2aa8
	13'h1555: q1 = 16'h48c1; // 0x2aaa
	13'h1556: q1 = 16'hd28e; // 0x2aac
	13'h1557: q1 = 16'h2241; // 0x2aae
	13'h1558: q1 = 16'h3229; // 0x2ab0
	13'h1559: q1 = 16'hfff4; // 0x2ab2
	13'h155a: q1 = 16'h1081; // 0x2ab4
	13'h155b: q1 = 16'h5245; // 0x2ab6
	13'h155c: q1 = 16'h60d4; // 0x2ab8
	13'h155d: q1 = 16'h4279; // 0x2aba
	13'h155e: q1 = 16'h0001; // 0x2abc
	13'h155f: q1 = 16'h7f20; // 0x2abe
	13'h1560: q1 = 16'h4a9f; // 0x2ac0
	13'h1561: q1 = 16'h4cdf; // 0x2ac2
	13'h1562: q1 = 16'h20f8; // 0x2ac4
	13'h1563: q1 = 16'h4e5e; // 0x2ac6
	13'h1564: q1 = 16'h4e75; // 0x2ac8
	13'h1565: q1 = 16'h4e56; // 0x2aca
	13'h1566: q1 = 16'hfffc; // 0x2acc
	13'h1567: q1 = 16'h536e; // 0x2ace
	13'h1568: q1 = 16'h0008; // 0x2ad0
	13'h1569: q1 = 16'h4a6e; // 0x2ad2
	13'h156a: q1 = 16'h0008; // 0x2ad4
	13'h156b: q1 = 16'h6740; // 0x2ad6
	13'h156c: q1 = 16'h4eb9; // 0x2ad8
	13'h156d: q1 = 16'h0000; // 0x2ada
	13'h156e: q1 = 16'h3fcc; // 0x2adc
	13'h156f: q1 = 16'h4eb9; // 0x2ade
	13'h1570: q1 = 16'h0000; // 0x2ae0
	13'h1571: q1 = 16'h909e; // 0x2ae2
	13'h1572: q1 = 16'h4eb9; // 0x2ae4
	13'h1573: q1 = 16'h0000; // 0x2ae6
	13'h1574: q1 = 16'h4820; // 0x2ae8
	13'h1575: q1 = 16'h4eb9; // 0x2aea
	13'h1576: q1 = 16'h0000; // 0x2aec
	13'h1577: q1 = 16'h18d0; // 0x2aee
	13'h1578: q1 = 16'h4eb9; // 0x2af0
	13'h1579: q1 = 16'h0000; // 0x2af2
	13'h157a: q1 = 16'h3434; // 0x2af4
	13'h157b: q1 = 16'h4ab9; // 0x2af6
	13'h157c: q1 = 16'h0001; // 0x2af8
	13'h157d: q1 = 16'h7fc2; // 0x2afa
	13'h157e: q1 = 16'h670e; // 0x2afc
	13'h157f: q1 = 16'h4a79; // 0x2afe
	13'h1580: q1 = 16'h0001; // 0x2b00
	13'h1581: q1 = 16'h7594; // 0x2b02
	13'h1582: q1 = 16'h6704; // 0x2b04
	13'h1583: q1 = 16'h7001; // 0x2b06
	13'h1584: q1 = 16'h601a; // 0x2b08
	13'h1585: q1 = 16'h60ea; // 0x2b0a
	13'h1586: q1 = 16'h23fc; // 0x2b0c
	13'h1587: q1 = 16'h0000; // 0x2b0e
	13'h1588: q1 = 16'h0002; // 0x2b10
	13'h1589: q1 = 16'h0001; // 0x2b12
	13'h158a: q1 = 16'h7fc2; // 0x2b14
	13'h158b: q1 = 16'h60b6; // 0x2b16
	13'h158c: q1 = 16'h23fc; // 0x2b18
	13'h158d: q1 = 16'h0000; // 0x2b1a
	13'h158e: q1 = 16'h0002; // 0x2b1c
	13'h158f: q1 = 16'h0001; // 0x2b1e
	13'h1590: q1 = 16'h7fc2; // 0x2b20
	13'h1591: q1 = 16'h4240; // 0x2b22
	13'h1592: q1 = 16'h4e5e; // 0x2b24
	13'h1593: q1 = 16'h4e75; // 0x2b26
	13'h1594: q1 = 16'h4e56; // 0x2b28
	13'h1595: q1 = 16'hffe0; // 0x2b2a
	13'h1596: q1 = 16'h48e7; // 0x2b2c
	13'h1597: q1 = 16'h0304; // 0x2b2e
	13'h1598: q1 = 16'h2a79; // 0x2b30
	13'h1599: q1 = 16'h0001; // 0x2b32
	13'h159a: q1 = 16'h7fb8; // 0x2b34
	13'h159b: q1 = 16'h0c55; // 0x2b36
	13'h159c: q1 = 16'h0005; // 0x2b38
	13'h159d: q1 = 16'h6d00; // 0x2b3a
	13'h159e: q1 = 16'h01bc; // 0x2b3c
	13'h159f: q1 = 16'h0c55; // 0x2b3e
	13'h15a0: q1 = 16'h0078; // 0x2b40
	13'h15a1: q1 = 16'h6e12; // 0x2b42
	13'h15a2: q1 = 16'h302d; // 0x2b44
	13'h15a3: q1 = 16'h0020; // 0x2b46
	13'h15a4: q1 = 16'h5a40; // 0x2b48
	13'h15a5: q1 = 16'hb055; // 0x2b4a
	13'h15a6: q1 = 16'h6f08; // 0x2b4c
	13'h15a7: q1 = 16'h4a6d; // 0x2b4e
	13'h15a8: q1 = 16'h0020; // 0x2b50
	13'h15a9: q1 = 16'h6e00; // 0x2b52
	13'h15aa: q1 = 16'h01a4; // 0x2b54
	13'h15ab: q1 = 16'h0c79; // 0x2b56
	13'h15ac: q1 = 16'h0018; // 0x2b58
	13'h15ad: q1 = 16'h0001; // 0x2b5a
	13'h15ae: q1 = 16'h81fc; // 0x2b5c
	13'h15af: q1 = 16'h6c00; // 0x2b5e
	13'h15b0: q1 = 16'h0198; // 0x2b60
	13'h15b1: q1 = 16'h0c79; // 0x2b62
	13'h15b2: q1 = 16'h0005; // 0x2b64
	13'h15b3: q1 = 16'h0001; // 0x2b66
	13'h15b4: q1 = 16'h7efc; // 0x2b68
	13'h15b5: q1 = 16'h6d00; // 0x2b6a
	13'h15b6: q1 = 16'h018c; // 0x2b6c
	13'h15b7: q1 = 16'h4a79; // 0x2b6e
	13'h15b8: q1 = 16'h0001; // 0x2b70
	13'h15b9: q1 = 16'h7f22; // 0x2b72
	13'h15ba: q1 = 16'h6700; // 0x2b74
	13'h15bb: q1 = 16'h0182; // 0x2b76
	13'h15bc: q1 = 16'h3b55; // 0x2b78
	13'h15bd: q1 = 16'h0020; // 0x2b7a
	13'h15be: q1 = 16'h4eb9; // 0x2b7c
	13'h15bf: q1 = 16'h0000; // 0x2b7e
	13'h15c0: q1 = 16'h0226; // 0x2b80
	13'h15c1: q1 = 16'h3ebc; // 0x2b82
	13'h15c2: q1 = 16'h0019; // 0x2b84
	13'h15c3: q1 = 16'h4eb9; // 0x2b86
	13'h15c4: q1 = 16'h0000; // 0x2b88
	13'h15c5: q1 = 16'h8a22; // 0x2b8a
	13'h15c6: q1 = 16'h7e2d; // 0x2b8c
	13'h15c7: q1 = 16'h23f9; // 0x2b8e
	13'h15c8: q1 = 16'h0000; // 0x2b90
	13'h15c9: q1 = 16'hce6c; // 0x2b92
	13'h15ca: q1 = 16'h0001; // 0x2b94
	13'h15cb: q1 = 16'h7f60; // 0x2b96
	13'h15cc: q1 = 16'h4ab9; // 0x2b98
	13'h15cd: q1 = 16'h0001; // 0x2b9a
	13'h15ce: q1 = 16'h7f60; // 0x2b9c
	13'h15cf: q1 = 16'h6756; // 0x2b9e
	13'h15d0: q1 = 16'h23fc; // 0x2ba0
	13'h15d1: q1 = 16'h0000; // 0x2ba2
	13'h15d2: q1 = 16'h0002; // 0x2ba4
	13'h15d3: q1 = 16'h0001; // 0x2ba6
	13'h15d4: q1 = 16'h7fc2; // 0x2ba8
	13'h15d5: q1 = 16'h3ebc; // 0x2baa
	13'h15d6: q1 = 16'h0035; // 0x2bac
	13'h15d7: q1 = 16'h200e; // 0x2bae
	13'h15d8: q1 = 16'hd0bc; // 0x2bb0
	13'h15d9: q1 = 16'hffff; // 0x2bb2
	13'h15da: q1 = 16'hffe0; // 0x2bb4
	13'h15db: q1 = 16'h2f00; // 0x2bb6
	13'h15dc: q1 = 16'h4eb9; // 0x2bb8
	13'h15dd: q1 = 16'h0000; // 0x2bba
	13'h15de: q1 = 16'h78f6; // 0x2bbc
	13'h15df: q1 = 16'h4a9f; // 0x2bbe
	13'h15e0: q1 = 16'h3e87; // 0x2bc0
	13'h15e1: q1 = 16'h4267; // 0x2bc2
	13'h15e2: q1 = 16'h3f3c; // 0x2bc4
	13'h15e3: q1 = 16'h0064; // 0x2bc6
	13'h15e4: q1 = 16'h3f3c; // 0x2bc8
	13'h15e5: q1 = 16'h0010; // 0x2bca
	13'h15e6: q1 = 16'h200e; // 0x2bcc
	13'h15e7: q1 = 16'hd0bc; // 0x2bce
	13'h15e8: q1 = 16'hffff; // 0x2bd0
	13'h15e9: q1 = 16'hffe0; // 0x2bd2
	13'h15ea: q1 = 16'h2f00; // 0x2bd4
	13'h15eb: q1 = 16'h4eb9; // 0x2bd6
	13'h15ec: q1 = 16'h0000; // 0x2bd8
	13'h15ed: q1 = 16'h026c; // 0x2bda
	13'h15ee: q1 = 16'hdefc; // 0x2bdc
	13'h15ef: q1 = 16'h000a; // 0x2bde
	13'h15f0: q1 = 16'h5247; // 0x2be0
	13'h15f1: q1 = 16'hbe7c; // 0x2be2
	13'h15f2: q1 = 16'h003f; // 0x2be4
	13'h15f3: q1 = 16'h6f02; // 0x2be6
	13'h15f4: q1 = 16'h7e2d; // 0x2be8
	13'h15f5: q1 = 16'h4ab9; // 0x2bea
	13'h15f6: q1 = 16'h0001; // 0x2bec
	13'h15f7: q1 = 16'h7fc2; // 0x2bee
	13'h15f8: q1 = 16'h6702; // 0x2bf0
	13'h15f9: q1 = 16'h60f6; // 0x2bf2
	13'h15fa: q1 = 16'h60a2; // 0x2bf4
	13'h15fb: q1 = 16'h33fc; // 0x2bf6
	13'h15fc: q1 = 16'h0001; // 0x2bf8
	13'h15fd: q1 = 16'h0001; // 0x2bfa
	13'h15fe: q1 = 16'h8676; // 0x2bfc
	13'h15ff: q1 = 16'h33f9; // 0x2bfe
	13'h1600: q1 = 16'h0001; // 0x2c00
	13'h1601: q1 = 16'h7eba; // 0x2c02
	13'h1602: q1 = 16'h0001; // 0x2c04
	13'h1603: q1 = 16'h8a76; // 0x2c06
	13'h1604: q1 = 16'h4eb9; // 0x2c08
	13'h1605: q1 = 16'h0000; // 0x2c0a
	13'h1606: q1 = 16'h0ea2; // 0x2c0c
	13'h1607: q1 = 16'h4eb9; // 0x2c0e
	13'h1608: q1 = 16'h0000; // 0x2c10
	13'h1609: q1 = 16'h41ae; // 0x2c12
	13'h160a: q1 = 16'h4eb9; // 0x2c14
	13'h160b: q1 = 16'h0000; // 0x2c16
	13'h160c: q1 = 16'hb3c6; // 0x2c18
	13'h160d: q1 = 16'h4eb9; // 0x2c1a
	13'h160e: q1 = 16'h0000; // 0x2c1c
	13'h160f: q1 = 16'h1e8a; // 0x2c1e
	13'h1610: q1 = 16'h4eb9; // 0x2c20
	13'h1611: q1 = 16'h0000; // 0x2c22
	13'h1612: q1 = 16'h4dee; // 0x2c24
	13'h1613: q1 = 16'h4eb9; // 0x2c26
	13'h1614: q1 = 16'h0000; // 0x2c28
	13'h1615: q1 = 16'h8330; // 0x2c2a
	13'h1616: q1 = 16'h4eb9; // 0x2c2c
	13'h1617: q1 = 16'h0000; // 0x2c2e
	13'h1618: q1 = 16'h5a9c; // 0x2c30
	13'h1619: q1 = 16'h4eb9; // 0x2c32
	13'h161a: q1 = 16'h0000; // 0x2c34
	13'h161b: q1 = 16'h2cba; // 0x2c36
	13'h161c: q1 = 16'h4eb9; // 0x2c38
	13'h161d: q1 = 16'h0000; // 0x2c3a
	13'h161e: q1 = 16'h90d4; // 0x2c3c
	13'h161f: q1 = 16'h33fc; // 0x2c3e
	13'h1620: q1 = 16'h0001; // 0x2c40
	13'h1621: q1 = 16'h0001; // 0x2c42
	13'h1622: q1 = 16'h7b9e; // 0x2c44
	13'h1623: q1 = 16'h33fc; // 0x2c46
	13'h1624: q1 = 16'h0001; // 0x2c48
	13'h1625: q1 = 16'h0001; // 0x2c4a
	13'h1626: q1 = 16'h86a8; // 0x2c4c
	13'h1627: q1 = 16'h4a79; // 0x2c4e
	13'h1628: q1 = 16'h0001; // 0x2c50
	13'h1629: q1 = 16'h86a8; // 0x2c52
	13'h162a: q1 = 16'h6722; // 0x2c54
	13'h162b: q1 = 16'h23fc; // 0x2c56
	13'h162c: q1 = 16'h0000; // 0x2c58
	13'h162d: q1 = 16'h0002; // 0x2c5a
	13'h162e: q1 = 16'h0001; // 0x2c5c
	13'h162f: q1 = 16'h7fc2; // 0x2c5e
	13'h1630: q1 = 16'h4eb9; // 0x2c60
	13'h1631: q1 = 16'h0000; // 0x2c62
	13'h1632: q1 = 16'h4820; // 0x2c64
	13'h1633: q1 = 16'h4eb9; // 0x2c66
	13'h1634: q1 = 16'h0000; // 0x2c68
	13'h1635: q1 = 16'h18d0; // 0x2c6a
	13'h1636: q1 = 16'h4ab9; // 0x2c6c
	13'h1637: q1 = 16'h0001; // 0x2c6e
	13'h1638: q1 = 16'h7fc2; // 0x2c70
	13'h1639: q1 = 16'h6702; // 0x2c72
	13'h163a: q1 = 16'h60f6; // 0x2c74
	13'h163b: q1 = 16'h60d6; // 0x2c76
	13'h163c: q1 = 16'h4279; // 0x2c78
	13'h163d: q1 = 16'h0001; // 0x2c7a
	13'h163e: q1 = 16'h7b9e; // 0x2c7c
	13'h163f: q1 = 16'h23fc; // 0x2c7e
	13'h1640: q1 = 16'h0000; // 0x2c80
	13'h1641: q1 = 16'h0002; // 0x2c82
	13'h1642: q1 = 16'h0001; // 0x2c84
	13'h1643: q1 = 16'h7fc2; // 0x2c86
	13'h1644: q1 = 16'h33fc; // 0x2c88
	13'h1645: q1 = 16'h0001; // 0x2c8a
	13'h1646: q1 = 16'h0001; // 0x2c8c
	13'h1647: q1 = 16'h805a; // 0x2c8e
	13'h1648: q1 = 16'h4eb9; // 0x2c90
	13'h1649: q1 = 16'h0000; // 0x2c92
	13'h164a: q1 = 16'h3434; // 0x2c94
	13'h164b: q1 = 16'h4eb9; // 0x2c96
	13'h164c: q1 = 16'h0000; // 0x2c98
	13'h164d: q1 = 16'h18d0; // 0x2c9a
	13'h164e: q1 = 16'h4eb9; // 0x2c9c
	13'h164f: q1 = 16'h0000; // 0x2c9e
	13'h1650: q1 = 16'h4820; // 0x2ca0
	13'h1651: q1 = 16'h4eb9; // 0x2ca2
	13'h1652: q1 = 16'h0000; // 0x2ca4
	13'h1653: q1 = 16'h909e; // 0x2ca6
	13'h1654: q1 = 16'h4eb9; // 0x2ca8
	13'h1655: q1 = 16'h0000; // 0x2caa
	13'h1656: q1 = 16'h3fcc; // 0x2cac
	13'h1657: q1 = 16'h4eb9; // 0x2cae
	13'h1658: q1 = 16'h0000; // 0x2cb0
	13'h1659: q1 = 16'h3396; // 0x2cb2
	13'h165a: q1 = 16'h4a40; // 0x2cb4
	13'h165b: q1 = 16'h6726; // 0x2cb6
	13'h165c: q1 = 16'h4eb9; // 0x2cb8
	13'h165d: q1 = 16'h0000; // 0x2cba
	13'h165e: q1 = 16'h4738; // 0x2cbc
	13'h165f: q1 = 16'h4a40; // 0x2cbe
	13'h1660: q1 = 16'h671c; // 0x2cc0
	13'h1661: q1 = 16'h4eb9; // 0x2cc2
	13'h1662: q1 = 16'h0000; // 0x2cc4
	13'h1663: q1 = 16'h16c2; // 0x2cc6
	13'h1664: q1 = 16'h4a40; // 0x2cc8
	13'h1665: q1 = 16'h6712; // 0x2cca
	13'h1666: q1 = 16'h4eb9; // 0x2ccc
	13'h1667: q1 = 16'h0000; // 0x2cce
	13'h1668: q1 = 16'h3fac; // 0x2cd0
	13'h1669: q1 = 16'h4a40; // 0x2cd2
	13'h166a: q1 = 16'h6708; // 0x2cd4
	13'h166b: q1 = 16'h4eb9; // 0x2cd6
	13'h166c: q1 = 16'h0000; // 0x2cd8
	13'h166d: q1 = 16'h18d0; // 0x2cda
	13'h166e: q1 = 16'h600c; // 0x2cdc
	13'h166f: q1 = 16'h4ab9; // 0x2cde
	13'h1670: q1 = 16'h0001; // 0x2ce0
	13'h1671: q1 = 16'h7fc2; // 0x2ce2
	13'h1672: q1 = 16'h6702; // 0x2ce4
	13'h1673: q1 = 16'h60f6; // 0x2ce6
	13'h1674: q1 = 16'h6094; // 0x2ce8
	13'h1675: q1 = 16'h4279; // 0x2cea
	13'h1676: q1 = 16'h0001; // 0x2cec
	13'h1677: q1 = 16'h8676; // 0x2cee
	13'h1678: q1 = 16'h33fc; // 0x2cf0
	13'h1679: q1 = 16'h0001; // 0x2cf2
	13'h167a: q1 = 16'h0001; // 0x2cf4
	13'h167b: q1 = 16'h7fc8; // 0x2cf6
	13'h167c: q1 = 16'h4a9f; // 0x2cf8
	13'h167d: q1 = 16'h4cdf; // 0x2cfa
	13'h167e: q1 = 16'h2080; // 0x2cfc
	13'h167f: q1 = 16'h4e5e; // 0x2cfe
	13'h1680: q1 = 16'h4e75; // 0x2d00
	13'h1681: q1 = 16'h4e56; // 0x2d02
	13'h1682: q1 = 16'hffb8; // 0x2d04
	13'h1683: q1 = 16'h48e7; // 0x2d06
	13'h1684: q1 = 16'h070c; // 0x2d08
	13'h1685: q1 = 16'h2a7c; // 0x2d0a
	13'h1686: q1 = 16'h0001; // 0x2d0c
	13'h1687: q1 = 16'h7f2c; // 0x2d0e
	13'h1688: q1 = 16'h33fc; // 0x2d10
	13'h1689: q1 = 16'h0001; // 0x2d12
	13'h168a: q1 = 16'h0001; // 0x2d14
	13'h168b: q1 = 16'h7faa; // 0x2d16
	13'h168c: q1 = 16'h4eb9; // 0x2d18
	13'h168d: q1 = 16'h0000; // 0x2d1a
	13'h168e: q1 = 16'h0226; // 0x2d1c
	13'h168f: q1 = 16'h2079; // 0x2d1e
	13'h1690: q1 = 16'h0001; // 0x2d20
	13'h1691: q1 = 16'h7fb8; // 0x2d22
	13'h1692: q1 = 16'h30bc; // 0x2d24
	13'h1693: q1 = 16'h0002; // 0x2d26
	13'h1694: q1 = 16'h2eb9; // 0x2d28
	13'h1695: q1 = 16'h0000; // 0x2d2a
	13'h1696: q1 = 16'hce70; // 0x2d2c
	13'h1697: q1 = 16'h4eb9; // 0x2d2e
	13'h1698: q1 = 16'h0000; // 0x2d30
	13'h1699: q1 = 16'h3a7c; // 0x2d32
	13'h169a: q1 = 16'h33f9; // 0x2d34
	13'h169b: q1 = 16'h0001; // 0x2d36
	13'h169c: q1 = 16'h8a76; // 0x2d38
	13'h169d: q1 = 16'h0001; // 0x2d3a
	13'h169e: q1 = 16'h7eba; // 0x2d3c
	13'h169f: q1 = 16'h33fc; // 0x2d3e
	13'h16a0: q1 = 16'hca43; // 0x2d40
	13'h16a1: q1 = 16'h0001; // 0x2d42
	13'h16a2: q1 = 16'h8a76; // 0x2d44
	13'h16a3: q1 = 16'h4eb9; // 0x2d46
	13'h16a4: q1 = 16'h0000; // 0x2d48
	13'h16a5: q1 = 16'h7aa4; // 0x2d4a
	13'h16a6: q1 = 16'h4a79; // 0x2d4c
	13'h16a7: q1 = 16'h0001; // 0x2d4e
	13'h16a8: q1 = 16'h7594; // 0x2d50
	13'h16a9: q1 = 16'h6600; // 0x2d52
	13'h16aa: q1 = 16'h06f4; // 0x2d54
	13'h16ab: q1 = 16'h4257; // 0x2d56
	13'h16ac: q1 = 16'h4eb9; // 0x2d58
	13'h16ad: q1 = 16'h0000; // 0x2d5a
	13'h16ae: q1 = 16'h5be0; // 0x2d5c
	13'h16af: q1 = 16'h4257; // 0x2d5e
	13'h16b0: q1 = 16'h4eb9; // 0x2d60
	13'h16b1: q1 = 16'h0000; // 0x2d62
	13'h16b2: q1 = 16'h8570; // 0x2d64
	13'h16b3: q1 = 16'h4257; // 0x2d66
	13'h16b4: q1 = 16'h4eb9; // 0x2d68
	13'h16b5: q1 = 16'h0000; // 0x2d6a
	13'h16b6: q1 = 16'h1710; // 0x2d6c
	13'h16b7: q1 = 16'h4257; // 0x2d6e
	13'h16b8: q1 = 16'h4eb9; // 0x2d70
	13'h16b9: q1 = 16'h0000; // 0x2d72
	13'h16ba: q1 = 16'h4770; // 0x2d74
	13'h16bb: q1 = 16'h4eb9; // 0x2d76
	13'h16bc: q1 = 16'h0000; // 0x2d78
	13'h16bd: q1 = 16'h42bc; // 0x2d7a
	13'h16be: q1 = 16'h3d7c; // 0x2d7c
	13'h16bf: q1 = 16'h0014; // 0x2d7e
	13'h16c0: q1 = 16'hfffe; // 0x2d80
	13'h16c1: q1 = 16'h7e01; // 0x2d82
	13'h16c2: q1 = 16'h3ebc; // 0x2d84
	13'h16c3: q1 = 16'h0005; // 0x2d86
	13'h16c4: q1 = 16'h4eb9; // 0x2d88
	13'h16c5: q1 = 16'h0000; // 0x2d8a
	13'h16c6: q1 = 16'h8a22; // 0x2d8c
	13'h16c7: q1 = 16'h23fc; // 0x2d8e
	13'h16c8: q1 = 16'h0000; // 0x2d90
	13'h16c9: q1 = 16'h0002; // 0x2d92
	13'h16ca: q1 = 16'h0001; // 0x2d94
	13'h16cb: q1 = 16'h7fc2; // 0x2d96
	13'h16cc: q1 = 16'h4eb9; // 0x2d98
	13'h16cd: q1 = 16'h0000; // 0x2d9a
	13'h16ce: q1 = 16'h18d0; // 0x2d9c
	13'h16cf: q1 = 16'h4eb9; // 0x2d9e
	13'h16d0: q1 = 16'h0000; // 0x2da0
	13'h16d1: q1 = 16'h2fb4; // 0x2da2
	13'h16d2: q1 = 16'h536e; // 0x2da4
	13'h16d3: q1 = 16'hfffe; // 0x2da6
	13'h16d4: q1 = 16'h4a6e; // 0x2da8
	13'h16d5: q1 = 16'hfffe; // 0x2daa
	13'h16d6: q1 = 16'h6600; // 0x2dac
	13'h16d7: q1 = 16'h00de; // 0x2dae
	13'h16d8: q1 = 16'hbe7c; // 0x2db0
	13'h16d9: q1 = 16'h0004; // 0x2db2
	13'h16da: q1 = 16'h6e00; // 0x2db4
	13'h16db: q1 = 16'h00f8; // 0x2db6
	13'h16dc: q1 = 16'h3e87; // 0x2db8
	13'h16dd: q1 = 16'h4eb9; // 0x2dba
	13'h16de: q1 = 16'h0000; // 0x2dbc
	13'h16df: q1 = 16'h1f1a; // 0x2dbe
	13'h16e0: q1 = 16'h3007; // 0x2dc0
	13'h16e1: q1 = 16'h6000; // 0x2dc2
	13'h16e2: q1 = 16'h0086; // 0x2dc4
	13'h16e3: q1 = 16'h2ebc; // 0x2dc6
	13'h16e4: q1 = 16'h0000; // 0x2dc8
	13'h16e5: q1 = 16'hce84; // 0x2dca
	13'h16e6: q1 = 16'h200e; // 0x2dcc
	13'h16e7: q1 = 16'hd0bc; // 0x2dce
	13'h16e8: q1 = 16'hffff; // 0x2dd0
	13'h16e9: q1 = 16'hffda; // 0x2dd2
	13'h16ea: q1 = 16'h2f00; // 0x2dd4
	13'h16eb: q1 = 16'h4eb9; // 0x2dd6
	13'h16ec: q1 = 16'h0000; // 0x2dd8
	13'h16ed: q1 = 16'h0750; // 0x2dda
	13'h16ee: q1 = 16'h4a9f; // 0x2ddc
	13'h16ef: q1 = 16'h3d7c; // 0x2dde
	13'h16f0: q1 = 16'h0015; // 0x2de0
	13'h16f1: q1 = 16'hfffc; // 0x2de2
	13'h16f2: q1 = 16'h6000; // 0x2de4
	13'h16f3: q1 = 16'h007a; // 0x2de6
	13'h16f4: q1 = 16'h2ebc; // 0x2de8
	13'h16f5: q1 = 16'h0000; // 0x2dea
	13'h16f6: q1 = 16'hce8a; // 0x2dec
	13'h16f7: q1 = 16'h200e; // 0x2dee
	13'h16f8: q1 = 16'hd0bc; // 0x2df0
	13'h16f9: q1 = 16'hffff; // 0x2df2
	13'h16fa: q1 = 16'hffda; // 0x2df4
	13'h16fb: q1 = 16'h2f00; // 0x2df6
	13'h16fc: q1 = 16'h4eb9; // 0x2df8
	13'h16fd: q1 = 16'h0000; // 0x2dfa
	13'h16fe: q1 = 16'h0750; // 0x2dfc
	13'h16ff: q1 = 16'h4a9f; // 0x2dfe
	13'h1700: q1 = 16'h3d7c; // 0x2e00
	13'h1701: q1 = 16'h0012; // 0x2e02
	13'h1702: q1 = 16'hfffc; // 0x2e04
	13'h1703: q1 = 16'h6058; // 0x2e06
	13'h1704: q1 = 16'h2ebc; // 0x2e08
	13'h1705: q1 = 16'h0000; // 0x2e0a
	13'h1706: q1 = 16'hce91; // 0x2e0c
	13'h1707: q1 = 16'h200e; // 0x2e0e
	13'h1708: q1 = 16'hd0bc; // 0x2e10
	13'h1709: q1 = 16'hffff; // 0x2e12
	13'h170a: q1 = 16'hffda; // 0x2e14
	13'h170b: q1 = 16'h2f00; // 0x2e16
	13'h170c: q1 = 16'h4eb9; // 0x2e18
	13'h170d: q1 = 16'h0000; // 0x2e1a
	13'h170e: q1 = 16'h0750; // 0x2e1c
	13'h170f: q1 = 16'h4a9f; // 0x2e1e
	13'h1710: q1 = 16'h3d7c; // 0x2e20
	13'h1711: q1 = 16'h000f; // 0x2e22
	13'h1712: q1 = 16'hfffc; // 0x2e24
	13'h1713: q1 = 16'h6038; // 0x2e26
	13'h1714: q1 = 16'h2ebc; // 0x2e28
	13'h1715: q1 = 16'h0000; // 0x2e2a
	13'h1716: q1 = 16'hce99; // 0x2e2c
	13'h1717: q1 = 16'h200e; // 0x2e2e
	13'h1718: q1 = 16'hd0bc; // 0x2e30
	13'h1719: q1 = 16'hffff; // 0x2e32
	13'h171a: q1 = 16'hffda; // 0x2e34
	13'h171b: q1 = 16'h2f00; // 0x2e36
	13'h171c: q1 = 16'h4eb9; // 0x2e38
	13'h171d: q1 = 16'h0000; // 0x2e3a
	13'h171e: q1 = 16'h0750; // 0x2e3c
	13'h171f: q1 = 16'h4a9f; // 0x2e3e
	13'h1720: q1 = 16'h3d7c; // 0x2e40
	13'h1721: q1 = 16'h000c; // 0x2e42
	13'h1722: q1 = 16'hfffc; // 0x2e44
	13'h1723: q1 = 16'h6018; // 0x2e46
	13'h1724: q1 = 16'h6016; // 0x2e48
	13'h1725: q1 = 16'h5340; // 0x2e4a
	13'h1726: q1 = 16'hb07c; // 0x2e4c
	13'h1727: q1 = 16'h0003; // 0x2e4e
	13'h1728: q1 = 16'h620e; // 0x2e50
	13'h1729: q1 = 16'he540; // 0x2e52
	13'h172a: q1 = 16'h3040; // 0x2e54
	13'h172b: q1 = 16'hd1fc; // 0x2e56
	13'h172c: q1 = 16'h0000; // 0x2e58
	13'h172d: q1 = 16'hce74; // 0x2e5a
	13'h172e: q1 = 16'h2050; // 0x2e5c
	13'h172f: q1 = 16'h4ed0; // 0x2e5e
	13'h1730: q1 = 16'h3ebc; // 0x2e60
	13'h1731: q1 = 16'h003e; // 0x2e62
	13'h1732: q1 = 16'h3f3c; // 0x2e64
	13'h1733: q1 = 16'h0007; // 0x2e66
	13'h1734: q1 = 16'h3f3c; // 0x2e68
	13'h1735: q1 = 16'h0005; // 0x2e6a
	13'h1736: q1 = 16'h3f2e; // 0x2e6c
	13'h1737: q1 = 16'hfffc; // 0x2e6e
	13'h1738: q1 = 16'h200e; // 0x2e70
	13'h1739: q1 = 16'hd0bc; // 0x2e72
	13'h173a: q1 = 16'hffff; // 0x2e74
	13'h173b: q1 = 16'hffda; // 0x2e76
	13'h173c: q1 = 16'h2f00; // 0x2e78
	13'h173d: q1 = 16'h4eb9; // 0x2e7a
	13'h173e: q1 = 16'h0000; // 0x2e7c
	13'h173f: q1 = 16'h026c; // 0x2e7e
	13'h1740: q1 = 16'hdefc; // 0x2e80
	13'h1741: q1 = 16'h000a; // 0x2e82
	13'h1742: q1 = 16'h5247; // 0x2e84
	13'h1743: q1 = 16'h3d7c; // 0x2e86
	13'h1744: q1 = 16'h0027; // 0x2e88
	13'h1745: q1 = 16'hfffe; // 0x2e8a
	13'h1746: q1 = 16'h4ab9; // 0x2e8c
	13'h1747: q1 = 16'h0001; // 0x2e8e
	13'h1748: q1 = 16'h7fc2; // 0x2e90
	13'h1749: q1 = 16'h670c; // 0x2e92
	13'h174a: q1 = 16'h4a79; // 0x2e94
	13'h174b: q1 = 16'h0001; // 0x2e96
	13'h174c: q1 = 16'h7594; // 0x2e98
	13'h174d: q1 = 16'h6600; // 0x2e9a
	13'h174e: q1 = 16'h05ac; // 0x2e9c
	13'h174f: q1 = 16'h60ec; // 0x2e9e
	13'h1750: q1 = 16'h23fc; // 0x2ea0
	13'h1751: q1 = 16'h0000; // 0x2ea2
	13'h1752: q1 = 16'h0002; // 0x2ea4
	13'h1753: q1 = 16'h0001; // 0x2ea6
	13'h1754: q1 = 16'h7fc2; // 0x2ea8
	13'h1755: q1 = 16'h6000; // 0x2eaa
	13'h1756: q1 = 16'hfeec; // 0x2eac
	13'h1757: q1 = 16'h33fc; // 0x2eae
	13'h1758: q1 = 16'h04d2; // 0x2eb0
	13'h1759: q1 = 16'h0001; // 0x2eb2
	13'h175a: q1 = 16'h8a76; // 0x2eb4
	13'h175b: q1 = 16'h3ebc; // 0x2eb6
	13'h175c: q1 = 16'h0015; // 0x2eb8
	13'h175d: q1 = 16'h4eb9; // 0x2eba
	13'h175e: q1 = 16'h0000; // 0x2ebc
	13'h175f: q1 = 16'h8a22; // 0x2ebe
	13'h1760: q1 = 16'h2079; // 0x2ec0
	13'h1761: q1 = 16'h0001; // 0x2ec2
	13'h1762: q1 = 16'h7fb8; // 0x2ec4
	13'h1763: q1 = 16'h30bc; // 0x2ec6
	13'h1764: q1 = 16'h0001; // 0x2ec8
	13'h1765: q1 = 16'h3ebc; // 0x2eca
	13'h1766: q1 = 16'h0001; // 0x2ecc
	13'h1767: q1 = 16'h4eb9; // 0x2ece
	13'h1768: q1 = 16'h0000; // 0x2ed0
	13'h1769: q1 = 16'h4770; // 0x2ed2
	13'h176a: q1 = 16'h4279; // 0x2ed4
	13'h176b: q1 = 16'h0001; // 0x2ed6
	13'h176c: q1 = 16'h8682; // 0x2ed8
	13'h176d: q1 = 16'h33fc; // 0x2eda
	13'h176e: q1 = 16'h0001; // 0x2edc
	13'h176f: q1 = 16'h0001; // 0x2ede
	13'h1770: q1 = 16'h8880; // 0x2ee0
	13'h1771: q1 = 16'h4279; // 0x2ee2
	13'h1772: q1 = 16'h0001; // 0x2ee4
	13'h1773: q1 = 16'h81fa; // 0x2ee6
	13'h1774: q1 = 16'h2ebc; // 0x2ee8
	13'h1775: q1 = 16'h0000; // 0x2eea
	13'h1776: q1 = 16'hce9f; // 0x2eec
	13'h1777: q1 = 16'h200e; // 0x2eee
	13'h1778: q1 = 16'hd0bc; // 0x2ef0
	13'h1779: q1 = 16'hffff; // 0x2ef2
	13'h177a: q1 = 16'hffda; // 0x2ef4
	13'h177b: q1 = 16'h2f00; // 0x2ef6
	13'h177c: q1 = 16'h4eb9; // 0x2ef8
	13'h177d: q1 = 16'h0000; // 0x2efa
	13'h177e: q1 = 16'h0750; // 0x2efc
	13'h177f: q1 = 16'h4a9f; // 0x2efe
	13'h1780: q1 = 16'h206d; // 0x2f00
	13'h1781: q1 = 16'h0024; // 0x2f02
	13'h1782: q1 = 16'h3010; // 0x2f04
	13'h1783: q1 = 16'h4281; // 0x2f06
	13'h1784: q1 = 16'h720a; // 0x2f08
	13'h1785: q1 = 16'he260; // 0x2f0a
	13'h1786: q1 = 16'h48c0; // 0x2f0c
	13'h1787: q1 = 16'hd08e; // 0x2f0e
	13'h1788: q1 = 16'h2040; // 0x2f10
	13'h1789: q1 = 16'h4a28; // 0x2f12
	13'h178a: q1 = 16'hffda; // 0x2f14
	13'h178b: q1 = 16'h6772; // 0x2f16
	13'h178c: q1 = 16'h4eb9; // 0x2f18
	13'h178d: q1 = 16'h0000; // 0x2f1a
	13'h178e: q1 = 16'h4820; // 0x2f1c
	13'h178f: q1 = 16'h4eb9; // 0x2f1e
	13'h1790: q1 = 16'h0000; // 0x2f20
	13'h1791: q1 = 16'h18d0; // 0x2f22
	13'h1792: q1 = 16'h4eb9; // 0x2f24
	13'h1793: q1 = 16'h0000; // 0x2f26
	13'h1794: q1 = 16'h2fb4; // 0x2f28
	13'h1795: q1 = 16'h206d; // 0x2f2a
	13'h1796: q1 = 16'h0024; // 0x2f2c
	13'h1797: q1 = 16'h3010; // 0x2f2e
	13'h1798: q1 = 16'h4281; // 0x2f30
	13'h1799: q1 = 16'h720a; // 0x2f32
	13'h179a: q1 = 16'he260; // 0x2f34
	13'h179b: q1 = 16'h6f30; // 0x2f36
	13'h179c: q1 = 16'h3ebc; // 0x2f38
	13'h179d: q1 = 16'h0031; // 0x2f3a
	13'h179e: q1 = 16'h206d; // 0x2f3c
	13'h179f: q1 = 16'h0024; // 0x2f3e
	13'h17a0: q1 = 16'h3010; // 0x2f40
	13'h17a1: q1 = 16'h4281; // 0x2f42
	13'h17a2: q1 = 16'h720a; // 0x2f44
	13'h17a3: q1 = 16'he260; // 0x2f46
	13'h17a4: q1 = 16'h48c0; // 0x2f48
	13'h17a5: q1 = 16'hd08e; // 0x2f4a
	13'h17a6: q1 = 16'h2040; // 0x2f4c
	13'h17a7: q1 = 16'h1028; // 0x2f4e
	13'h17a8: q1 = 16'hffda; // 0x2f50
	13'h17a9: q1 = 16'h4880; // 0x2f52
	13'h17aa: q1 = 16'h3f00; // 0x2f54
	13'h17ab: q1 = 16'h3f3c; // 0x2f56
	13'h17ac: q1 = 16'h1c00; // 0x2f58
	13'h17ad: q1 = 16'h206d; // 0x2f5a
	13'h17ae: q1 = 16'h0024; // 0x2f5c
	13'h17af: q1 = 16'h3f10; // 0x2f5e
	13'h17b0: q1 = 16'h4eb9; // 0x2f60
	13'h17b1: q1 = 16'h0000; // 0x2f62
	13'h17b2: q1 = 16'h3f80; // 0x2f64
	13'h17b3: q1 = 16'h5c4f; // 0x2f66
	13'h17b4: q1 = 16'h4ab9; // 0x2f68
	13'h17b5: q1 = 16'h0001; // 0x2f6a
	13'h17b6: q1 = 16'h7fc2; // 0x2f6c
	13'h17b7: q1 = 16'h670c; // 0x2f6e
	13'h17b8: q1 = 16'h4a79; // 0x2f70
	13'h17b9: q1 = 16'h0001; // 0x2f72
	13'h17ba: q1 = 16'h7594; // 0x2f74
	13'h17bb: q1 = 16'h6600; // 0x2f76
	13'h17bc: q1 = 16'h04d0; // 0x2f78
	13'h17bd: q1 = 16'h60ec; // 0x2f7a
	13'h17be: q1 = 16'h23fc; // 0x2f7c
	13'h17bf: q1 = 16'h0000; // 0x2f7e
	13'h17c0: q1 = 16'h0002; // 0x2f80
	13'h17c1: q1 = 16'h0001; // 0x2f82
	13'h17c2: q1 = 16'h7fc2; // 0x2f84
	13'h17c3: q1 = 16'h6000; // 0x2f86
	13'h17c4: q1 = 16'hff78; // 0x2f88
	13'h17c5: q1 = 16'h3d7c; // 0x2f8a
	13'h17c6: q1 = 16'h0028; // 0x2f8c
	13'h17c7: q1 = 16'hfffe; // 0x2f8e
	13'h17c8: q1 = 16'h536e; // 0x2f90
	13'h17c9: q1 = 16'hfffe; // 0x2f92
	13'h17ca: q1 = 16'h4a6e; // 0x2f94
	13'h17cb: q1 = 16'hfffe; // 0x2f96
	13'h17cc: q1 = 16'h6748; // 0x2f98
	13'h17cd: q1 = 16'h4279; // 0x2f9a
	13'h17ce: q1 = 16'h0001; // 0x2f9c
	13'h17cf: q1 = 16'h8880; // 0x2f9e
	13'h17d0: q1 = 16'h0c79; // 0x2fa0
	13'h17d1: q1 = 16'h0024; // 0x2fa2
	13'h17d2: q1 = 16'h0001; // 0x2fa4
	13'h17d3: q1 = 16'h8682; // 0x2fa6
	13'h17d4: q1 = 16'h6c06; // 0x2fa8
	13'h17d5: q1 = 16'h5279; // 0x2faa
	13'h17d6: q1 = 16'h0001; // 0x2fac
	13'h17d7: q1 = 16'h8682; // 0x2fae
	13'h17d8: q1 = 16'h4eb9; // 0x2fb0
	13'h17d9: q1 = 16'h0000; // 0x2fb2
	13'h17da: q1 = 16'h4820; // 0x2fb4
	13'h17db: q1 = 16'h4eb9; // 0x2fb6
	13'h17dc: q1 = 16'h0000; // 0x2fb8
	13'h17dd: q1 = 16'h18d0; // 0x2fba
	13'h17de: q1 = 16'h4eb9; // 0x2fbc
	13'h17df: q1 = 16'h0000; // 0x2fbe
	13'h17e0: q1 = 16'h2fb4; // 0x2fc0
	13'h17e1: q1 = 16'h4ab9; // 0x2fc2
	13'h17e2: q1 = 16'h0001; // 0x2fc4
	13'h17e3: q1 = 16'h7fc2; // 0x2fc6
	13'h17e4: q1 = 16'h670c; // 0x2fc8
	13'h17e5: q1 = 16'h4a79; // 0x2fca
	13'h17e6: q1 = 16'h0001; // 0x2fcc
	13'h17e7: q1 = 16'h7594; // 0x2fce
	13'h17e8: q1 = 16'h6600; // 0x2fd0
	13'h17e9: q1 = 16'h0476; // 0x2fd2
	13'h17ea: q1 = 16'h60ec; // 0x2fd4
	13'h17eb: q1 = 16'h23fc; // 0x2fd6
	13'h17ec: q1 = 16'h0000; // 0x2fd8
	13'h17ed: q1 = 16'h0002; // 0x2fda
	13'h17ee: q1 = 16'h0001; // 0x2fdc
	13'h17ef: q1 = 16'h7fc2; // 0x2fde
	13'h17f0: q1 = 16'h60ae; // 0x2fe0
	13'h17f1: q1 = 16'h33fc; // 0x2fe2
	13'h17f2: q1 = 16'h0001; // 0x2fe4
	13'h17f3: q1 = 16'h0001; // 0x2fe6
	13'h17f4: q1 = 16'h806e; // 0x2fe8
	13'h17f5: q1 = 16'h3ebc; // 0x2fea
	13'h17f6: q1 = 16'h0002; // 0x2fec
	13'h17f7: q1 = 16'h4eb9; // 0x2fee
	13'h17f8: q1 = 16'h0000; // 0x2ff0
	13'h17f9: q1 = 16'h5be0; // 0x2ff2
	13'h17fa: q1 = 16'h3ebc; // 0x2ff4
	13'h17fb: q1 = 16'h0002; // 0x2ff6
	13'h17fc: q1 = 16'h4eb9; // 0x2ff8
	13'h17fd: q1 = 16'h0000; // 0x2ffa
	13'h17fe: q1 = 16'h1710; // 0x2ffc
	13'h17ff: q1 = 16'h4eb9; // 0x2ffe
	13'h1800: q1 = 16'h0000; // 0x3000
	13'h1801: q1 = 16'h2fb4; // 0x3002
	13'h1802: q1 = 16'h4eb9; // 0x3004
	13'h1803: q1 = 16'h0000; // 0x3006
	13'h1804: q1 = 16'h4820; // 0x3008
	13'h1805: q1 = 16'h4eb9; // 0x300a
	13'h1806: q1 = 16'h0000; // 0x300c
	13'h1807: q1 = 16'h18d0; // 0x300e
	13'h1808: q1 = 16'h3ebc; // 0x3010
	13'h1809: q1 = 16'h0018; // 0x3012
	13'h180a: q1 = 16'h3f3c; // 0x3014
	13'h180b: q1 = 16'h0004; // 0x3016
	13'h180c: q1 = 16'h4eb9; // 0x3018
	13'h180d: q1 = 16'h0000; // 0x301a
	13'h180e: q1 = 16'h01e4; // 0x301c
	13'h180f: q1 = 16'h4a5f; // 0x301e
	13'h1810: q1 = 16'h3ebc; // 0x3020
	13'h1811: q1 = 16'h0016; // 0x3022
	13'h1812: q1 = 16'h4eb9; // 0x3024
	13'h1813: q1 = 16'h0000; // 0x3026
	13'h1814: q1 = 16'h8a22; // 0x3028
	13'h1815: q1 = 16'h4ab9; // 0x302a
	13'h1816: q1 = 16'h0001; // 0x302c
	13'h1817: q1 = 16'h7fc2; // 0x302e
	13'h1818: q1 = 16'h670c; // 0x3030
	13'h1819: q1 = 16'h4a79; // 0x3032
	13'h181a: q1 = 16'h0001; // 0x3034
	13'h181b: q1 = 16'h7594; // 0x3036
	13'h181c: q1 = 16'h6600; // 0x3038
	13'h181d: q1 = 16'h040e; // 0x303a
	13'h181e: q1 = 16'h60ec; // 0x303c
	13'h181f: q1 = 16'h3d7c; // 0x303e
	13'h1820: q1 = 16'h003c; // 0x3040
	13'h1821: q1 = 16'hfffe; // 0x3042
	13'h1822: q1 = 16'h536e; // 0x3044
	13'h1823: q1 = 16'hfffe; // 0x3046
	13'h1824: q1 = 16'h4a6e; // 0x3048
	13'h1825: q1 = 16'hfffe; // 0x304a
	13'h1826: q1 = 16'h6732; // 0x304c
	13'h1827: q1 = 16'h4eb9; // 0x304e
	13'h1828: q1 = 16'h0000; // 0x3050
	13'h1829: q1 = 16'h4820; // 0x3052
	13'h182a: q1 = 16'h4eb9; // 0x3054
	13'h182b: q1 = 16'h0000; // 0x3056
	13'h182c: q1 = 16'h18d0; // 0x3058
	13'h182d: q1 = 16'h4eb9; // 0x305a
	13'h182e: q1 = 16'h0000; // 0x305c
	13'h182f: q1 = 16'h2fb4; // 0x305e
	13'h1830: q1 = 16'h4ab9; // 0x3060
	13'h1831: q1 = 16'h0001; // 0x3062
	13'h1832: q1 = 16'h7fc2; // 0x3064
	13'h1833: q1 = 16'h670c; // 0x3066
	13'h1834: q1 = 16'h4a79; // 0x3068
	13'h1835: q1 = 16'h0001; // 0x306a
	13'h1836: q1 = 16'h7594; // 0x306c
	13'h1837: q1 = 16'h6600; // 0x306e
	13'h1838: q1 = 16'h03d8; // 0x3070
	13'h1839: q1 = 16'h60ec; // 0x3072
	13'h183a: q1 = 16'h23fc; // 0x3074
	13'h183b: q1 = 16'h0000; // 0x3076
	13'h183c: q1 = 16'h0002; // 0x3078
	13'h183d: q1 = 16'h0001; // 0x307a
	13'h183e: q1 = 16'h7fc2; // 0x307c
	13'h183f: q1 = 16'h60c4; // 0x307e
	13'h1840: q1 = 16'h4eb9; // 0x3080
	13'h1841: q1 = 16'h0000; // 0x3082
	13'h1842: q1 = 16'h41ae; // 0x3084
	13'h1843: q1 = 16'h4eb9; // 0x3086
	13'h1844: q1 = 16'h0000; // 0x3088
	13'h1845: q1 = 16'h90d4; // 0x308a
	13'h1846: q1 = 16'h7c06; // 0x308c
	13'h1847: q1 = 16'hbc7c; // 0x308e
	13'h1848: q1 = 16'h0009; // 0x3090
	13'h1849: q1 = 16'h6e0c; // 0x3092
	13'h184a: q1 = 16'h3e86; // 0x3094
	13'h184b: q1 = 16'h4eb9; // 0x3096
	13'h184c: q1 = 16'h0000; // 0x3098
	13'h184d: q1 = 16'h8a22; // 0x309a
	13'h184e: q1 = 16'h5246; // 0x309c
	13'h184f: q1 = 16'h60ee; // 0x309e
	13'h1850: q1 = 16'h3ebc; // 0x30a0
	13'h1851: q1 = 16'h0096; // 0x30a2
	13'h1852: q1 = 16'h4eb9; // 0x30a4
	13'h1853: q1 = 16'h0000; // 0x30a6
	13'h1854: q1 = 16'h6aca; // 0x30a8
	13'h1855: q1 = 16'h4a40; // 0x30aa
	13'h1856: q1 = 16'h6600; // 0x30ac
	13'h1857: q1 = 16'h039a; // 0x30ae
	13'h1858: q1 = 16'h3ebc; // 0x30b0
	13'h1859: q1 = 16'h0007; // 0x30b2
	13'h185a: q1 = 16'h3f3c; // 0x30b4
	13'h185b: q1 = 16'h0004; // 0x30b6
	13'h185c: q1 = 16'h4eb9; // 0x30b8
	13'h185d: q1 = 16'h0000; // 0x30ba
	13'h185e: q1 = 16'h01e4; // 0x30bc
	13'h185f: q1 = 16'h4a5f; // 0x30be
	13'h1860: q1 = 16'h3ebc; // 0x30c0
	13'h1861: q1 = 16'h0003; // 0x30c2
	13'h1862: q1 = 16'h4eb9; // 0x30c4
	13'h1863: q1 = 16'h0000; // 0x30c6
	13'h1864: q1 = 16'h8570; // 0x30c8
	13'h1865: q1 = 16'h3ebc; // 0x30ca
	13'h1866: q1 = 16'h0003; // 0x30cc
	13'h1867: q1 = 16'h4eb9; // 0x30ce
	13'h1868: q1 = 16'h0000; // 0x30d0
	13'h1869: q1 = 16'h5be0; // 0x30d2
	13'h186a: q1 = 16'h3ebc; // 0x30d4
	13'h186b: q1 = 16'h005a; // 0x30d6
	13'h186c: q1 = 16'h4eb9; // 0x30d8
	13'h186d: q1 = 16'h0000; // 0x30da
	13'h186e: q1 = 16'h6aca; // 0x30dc
	13'h186f: q1 = 16'h4a40; // 0x30de
	13'h1870: q1 = 16'h6600; // 0x30e0
	13'h1871: q1 = 16'h0366; // 0x30e2
	13'h1872: q1 = 16'h3ebc; // 0x30e4
	13'h1873: q1 = 16'h0004; // 0x30e6
	13'h1874: q1 = 16'h4eb9; // 0x30e8
	13'h1875: q1 = 16'h0000; // 0x30ea
	13'h1876: q1 = 16'h8570; // 0x30ec
	13'h1877: q1 = 16'h7c0a; // 0x30ee
	13'h1878: q1 = 16'hbc7c; // 0x30f0
	13'h1879: q1 = 16'h000c; // 0x30f2
	13'h187a: q1 = 16'h6e0c; // 0x30f4
	13'h187b: q1 = 16'h3e86; // 0x30f6
	13'h187c: q1 = 16'h4eb9; // 0x30f8
	13'h187d: q1 = 16'h0000; // 0x30fa
	13'h187e: q1 = 16'h8a22; // 0x30fc
	13'h187f: q1 = 16'h5246; // 0x30fe
	13'h1880: q1 = 16'h60ee; // 0x3100
	13'h1881: q1 = 16'h3ebc; // 0x3102
	13'h1882: q1 = 16'h005a; // 0x3104
	13'h1883: q1 = 16'h4eb9; // 0x3106
	13'h1884: q1 = 16'h0000; // 0x3108
	13'h1885: q1 = 16'h6aca; // 0x310a
	13'h1886: q1 = 16'h4a40; // 0x310c
	13'h1887: q1 = 16'h6600; // 0x310e
	13'h1888: q1 = 16'h0338; // 0x3110
	13'h1889: q1 = 16'h3ebc; // 0x3112
	13'h188a: q1 = 16'h0007; // 0x3114
	13'h188b: q1 = 16'h3f3c; // 0x3116
	13'h188c: q1 = 16'h0007; // 0x3118
	13'h188d: q1 = 16'h4eb9; // 0x311a
	13'h188e: q1 = 16'h0000; // 0x311c
	13'h188f: q1 = 16'h01e4; // 0x311e
	13'h1890: q1 = 16'h4a5f; // 0x3120
	13'h1891: q1 = 16'h3ebc; // 0x3122
	13'h1892: q1 = 16'h000d; // 0x3124
	13'h1893: q1 = 16'h4eb9; // 0x3126
	13'h1894: q1 = 16'h0000; // 0x3128
	13'h1895: q1 = 16'h8a22; // 0x312a
	13'h1896: q1 = 16'h3ebc; // 0x312c
	13'h1897: q1 = 16'h000e; // 0x312e
	13'h1898: q1 = 16'h4eb9; // 0x3130
	13'h1899: q1 = 16'h0000; // 0x3132
	13'h189a: q1 = 16'h8a22; // 0x3134
	13'h189b: q1 = 16'h3ebc; // 0x3136
	13'h189c: q1 = 16'h0078; // 0x3138
	13'h189d: q1 = 16'h4eb9; // 0x313a
	13'h189e: q1 = 16'h0000; // 0x313c
	13'h189f: q1 = 16'h6aca; // 0x313e
	13'h18a0: q1 = 16'h4a40; // 0x3140
	13'h18a1: q1 = 16'h6600; // 0x3142
	13'h18a2: q1 = 16'h0304; // 0x3144
	13'h18a3: q1 = 16'h2079; // 0x3146
	13'h18a4: q1 = 16'h0001; // 0x3148
	13'h18a5: q1 = 16'h7fb8; // 0x314a
	13'h18a6: q1 = 16'h30bc; // 0x314c
	13'h18a7: q1 = 16'h0002; // 0x314e
	13'h18a8: q1 = 16'h3ebc; // 0x3150
	13'h18a9: q1 = 16'h0005; // 0x3152
	13'h18aa: q1 = 16'h4eb9; // 0x3154
	13'h18ab: q1 = 16'h0000; // 0x3156
	13'h18ac: q1 = 16'h1710; // 0x3158
	13'h18ad: q1 = 16'h3ebc; // 0x315a
	13'h18ae: q1 = 16'h000f; // 0x315c
	13'h18af: q1 = 16'h4eb9; // 0x315e
	13'h18b0: q1 = 16'h0000; // 0x3160
	13'h18b1: q1 = 16'h8a22; // 0x3162
	13'h18b2: q1 = 16'h3ebc; // 0x3164
	13'h18b3: q1 = 16'h0010; // 0x3166
	13'h18b4: q1 = 16'h4eb9; // 0x3168
	13'h18b5: q1 = 16'h0000; // 0x316a
	13'h18b6: q1 = 16'h8a22; // 0x316c
	13'h18b7: q1 = 16'h3ebc; // 0x316e
	13'h18b8: q1 = 16'h0078; // 0x3170
	13'h18b9: q1 = 16'h4eb9; // 0x3172
	13'h18ba: q1 = 16'h0000; // 0x3174
	13'h18bb: q1 = 16'h6aca; // 0x3176
	13'h18bc: q1 = 16'h4a40; // 0x3178
	13'h18bd: q1 = 16'h6600; // 0x317a
	13'h18be: q1 = 16'h02cc; // 0x317c
	13'h18bf: q1 = 16'h3ebc; // 0x317e
	13'h18c0: q1 = 16'h0011; // 0x3180
	13'h18c1: q1 = 16'h4eb9; // 0x3182
	13'h18c2: q1 = 16'h0000; // 0x3184
	13'h18c3: q1 = 16'h8a22; // 0x3186
	13'h18c4: q1 = 16'h3ebc; // 0x3188
	13'h18c5: q1 = 16'h0012; // 0x318a
	13'h18c6: q1 = 16'h4eb9; // 0x318c
	13'h18c7: q1 = 16'h0000; // 0x318e
	13'h18c8: q1 = 16'h8a22; // 0x3190
	13'h18c9: q1 = 16'h3ebc; // 0x3192
	13'h18ca: q1 = 16'h0005; // 0x3194
	13'h18cb: q1 = 16'h3f3c; // 0x3196
	13'h18cc: q1 = 16'h0005; // 0x3198
	13'h18cd: q1 = 16'h4eb9; // 0x319a
	13'h18ce: q1 = 16'h0000; // 0x319c
	13'h18cf: q1 = 16'h01e4; // 0x319e
	13'h18d0: q1 = 16'h4a5f; // 0x31a0
	13'h18d1: q1 = 16'h3ebc; // 0x31a2
	13'h18d2: q1 = 16'h005a; // 0x31a4
	13'h18d3: q1 = 16'h4eb9; // 0x31a6
	13'h18d4: q1 = 16'h0000; // 0x31a8
	13'h18d5: q1 = 16'h6aca; // 0x31aa
	13'h18d6: q1 = 16'h4a40; // 0x31ac
	13'h18d7: q1 = 16'h6600; // 0x31ae
	13'h18d8: q1 = 16'h0298; // 0x31b0
	13'h18d9: q1 = 16'h3ebc; // 0x31b2
	13'h18da: q1 = 16'h0013; // 0x31b4
	13'h18db: q1 = 16'h4eb9; // 0x31b6
	13'h18dc: q1 = 16'h0000; // 0x31b8
	13'h18dd: q1 = 16'h8a22; // 0x31ba
	13'h18de: q1 = 16'h3ebc; // 0x31bc
	13'h18df: q1 = 16'h0014; // 0x31be
	13'h18e0: q1 = 16'h4eb9; // 0x31c0
	13'h18e1: q1 = 16'h0000; // 0x31c2
	13'h18e2: q1 = 16'h8a22; // 0x31c4
	13'h18e3: q1 = 16'h3ebc; // 0x31c6
	13'h18e4: q1 = 16'h0006; // 0x31c8
	13'h18e5: q1 = 16'h4eb9; // 0x31ca
	13'h18e6: q1 = 16'h0000; // 0x31cc
	13'h18e7: q1 = 16'h5be0; // 0x31ce
	13'h18e8: q1 = 16'h3ebc; // 0x31d0
	13'h18e9: q1 = 16'h005a; // 0x31d2
	13'h18ea: q1 = 16'h4eb9; // 0x31d4
	13'h18eb: q1 = 16'h0000; // 0x31d6
	13'h18ec: q1 = 16'h6aca; // 0x31d8
	13'h18ed: q1 = 16'h4a40; // 0x31da
	13'h18ee: q1 = 16'h6600; // 0x31dc
	13'h18ef: q1 = 16'h026a; // 0x31de
	13'h18f0: q1 = 16'h3ebc; // 0x31e0
	13'h18f1: q1 = 16'h0007; // 0x31e2
	13'h18f2: q1 = 16'h3f3c; // 0x31e4
	13'h18f3: q1 = 16'h0004; // 0x31e6
	13'h18f4: q1 = 16'h4eb9; // 0x31e8
	13'h18f5: q1 = 16'h0000; // 0x31ea
	13'h18f6: q1 = 16'h01e4; // 0x31ec
	13'h18f7: q1 = 16'h4a5f; // 0x31ee
	13'h18f8: q1 = 16'h3ebc; // 0x31f0
	13'h18f9: q1 = 16'h0005; // 0x31f2
	13'h18fa: q1 = 16'h4eb9; // 0x31f4
	13'h18fb: q1 = 16'h0000; // 0x31f6
	13'h18fc: q1 = 16'h1710; // 0x31f8
	13'h18fd: q1 = 16'h3039; // 0x31fa
	13'h18fe: q1 = 16'h0001; // 0x31fc
	13'h18ff: q1 = 16'h7580; // 0x31fe
	13'h1900: q1 = 16'hd079; // 0x3200
	13'h1901: q1 = 16'h0001; // 0x3202
	13'h1902: q1 = 16'h7582; // 0x3204
	13'h1903: q1 = 16'hd079; // 0x3206
	13'h1904: q1 = 16'h0001; // 0x3208
	13'h1905: q1 = 16'h7586; // 0x320a
	13'h1906: q1 = 16'h6f0a; // 0x320c
	13'h1907: q1 = 16'h3ebc; // 0x320e
	13'h1908: q1 = 16'h0004; // 0x3210
	13'h1909: q1 = 16'h4eb9; // 0x3212
	13'h190a: q1 = 16'h0000; // 0x3214
	13'h190b: q1 = 16'h8a22; // 0x3216
	13'h190c: q1 = 16'h7c06; // 0x3218
	13'h190d: q1 = 16'h4a79; // 0x321a
	13'h190e: q1 = 16'h0001; // 0x321c
	13'h190f: q1 = 16'h7580; // 0x321e
	13'h1910: q1 = 16'h6f00; // 0x3220
	13'h1911: q1 = 16'h00d6; // 0x3222
	13'h1912: q1 = 16'h3ebc; // 0x3224
	13'h1913: q1 = 16'h0010; // 0x3226
	13'h1914: q1 = 16'h200e; // 0x3228
	13'h1915: q1 = 16'hd0bc; // 0x322a
	13'h1916: q1 = 16'hffff; // 0x322c
	13'h1917: q1 = 16'hffda; // 0x322e
	13'h1918: q1 = 16'h2f00; // 0x3230
	13'h1919: q1 = 16'h4eb9; // 0x3232
	13'h191a: q1 = 16'h0000; // 0x3234
	13'h191b: q1 = 16'h78f6; // 0x3236
	13'h191c: q1 = 16'h4a9f; // 0x3238
	13'h191d: q1 = 16'h200e; // 0x323a
	13'h191e: q1 = 16'hd0bc; // 0x323c
	13'h191f: q1 = 16'hffff; // 0x323e
	13'h1920: q1 = 16'hffda; // 0x3240
	13'h1921: q1 = 16'h2e80; // 0x3242
	13'h1922: q1 = 16'h3f39; // 0x3244
	13'h1923: q1 = 16'h0001; // 0x3246
	13'h1924: q1 = 16'h7580; // 0x3248
	13'h1925: q1 = 16'h4eb9; // 0x324a
	13'h1926: q1 = 16'h0000; // 0x324c
	13'h1927: q1 = 16'h0798; // 0x324e
	13'h1928: q1 = 16'h4a5f; // 0x3250
	13'h1929: q1 = 16'h3ebc; // 0x3252
	13'h192a: q1 = 16'h0011; // 0x3254
	13'h192b: q1 = 16'h200e; // 0x3256
	13'h192c: q1 = 16'hd0bc; // 0x3258
	13'h192d: q1 = 16'hffff; // 0x325a
	13'h192e: q1 = 16'hffb8; // 0x325c
	13'h192f: q1 = 16'h2f00; // 0x325e
	13'h1930: q1 = 16'h4eb9; // 0x3260
	13'h1931: q1 = 16'h0000; // 0x3262
	13'h1932: q1 = 16'h78f6; // 0x3264
	13'h1933: q1 = 16'h4a9f; // 0x3266
	13'h1934: q1 = 16'h200e; // 0x3268
	13'h1935: q1 = 16'hd0bc; // 0x326a
	13'h1936: q1 = 16'hffff; // 0x326c
	13'h1937: q1 = 16'hffb8; // 0x326e
	13'h1938: q1 = 16'h2e80; // 0x3270
	13'h1939: q1 = 16'h200e; // 0x3272
	13'h193a: q1 = 16'hd0bc; // 0x3274
	13'h193b: q1 = 16'hffff; // 0x3276
	13'h193c: q1 = 16'hffda; // 0x3278
	13'h193d: q1 = 16'h2f00; // 0x327a
	13'h193e: q1 = 16'h4eb9; // 0x327c
	13'h193f: q1 = 16'h0000; // 0x327e
	13'h1940: q1 = 16'h0770; // 0x3280
	13'h1941: q1 = 16'h4a9f; // 0x3282
	13'h1942: q1 = 16'h3039; // 0x3284
	13'h1943: q1 = 16'h0001; // 0x3286
	13'h1944: q1 = 16'h7582; // 0x3288
	13'h1945: q1 = 16'hd079; // 0x328a
	13'h1946: q1 = 16'h0001; // 0x328c
	13'h1947: q1 = 16'h7586; // 0x328e
	13'h1948: q1 = 16'h6f42; // 0x3290
	13'h1949: q1 = 16'h4a79; // 0x3292
	13'h194a: q1 = 16'h0001; // 0x3294
	13'h194b: q1 = 16'h7582; // 0x3296
	13'h194c: q1 = 16'h6708; // 0x3298
	13'h194d: q1 = 16'h4a79; // 0x329a
	13'h194e: q1 = 16'h0001; // 0x329c
	13'h194f: q1 = 16'h7586; // 0x329e
	13'h1950: q1 = 16'h6632; // 0x32a0
	13'h1951: q1 = 16'h3ebc; // 0x32a2
	13'h1952: q1 = 16'h0012; // 0x32a4
	13'h1953: q1 = 16'h200e; // 0x32a6
	13'h1954: q1 = 16'hd0bc; // 0x32a8
	13'h1955: q1 = 16'hffff; // 0x32aa
	13'h1956: q1 = 16'hffb8; // 0x32ac
	13'h1957: q1 = 16'h2f00; // 0x32ae
	13'h1958: q1 = 16'h4eb9; // 0x32b0
	13'h1959: q1 = 16'h0000; // 0x32b2
	13'h195a: q1 = 16'h78f6; // 0x32b4
	13'h195b: q1 = 16'h4a9f; // 0x32b6
	13'h195c: q1 = 16'h200e; // 0x32b8
	13'h195d: q1 = 16'hd0bc; // 0x32ba
	13'h195e: q1 = 16'hffff; // 0x32bc
	13'h195f: q1 = 16'hffb8; // 0x32be
	13'h1960: q1 = 16'h2e80; // 0x32c0
	13'h1961: q1 = 16'h200e; // 0x32c2
	13'h1962: q1 = 16'hd0bc; // 0x32c4
	13'h1963: q1 = 16'hffff; // 0x32c6
	13'h1964: q1 = 16'hffda; // 0x32c8
	13'h1965: q1 = 16'h2f00; // 0x32ca
	13'h1966: q1 = 16'h4eb9; // 0x32cc
	13'h1967: q1 = 16'h0000; // 0x32ce
	13'h1968: q1 = 16'h0770; // 0x32d0
	13'h1969: q1 = 16'h4a9f; // 0x32d2
	13'h196a: q1 = 16'h3ebc; // 0x32d4
	13'h196b: q1 = 16'h0032; // 0x32d6
	13'h196c: q1 = 16'h3f3c; // 0x32d8
	13'h196d: q1 = 16'h0020; // 0x32da
	13'h196e: q1 = 16'h3f3c; // 0x32dc
	13'h196f: q1 = 16'h0064; // 0x32de
	13'h1970: q1 = 16'h3f06; // 0x32e0
	13'h1971: q1 = 16'h5346; // 0x32e2
	13'h1972: q1 = 16'h200e; // 0x32e4
	13'h1973: q1 = 16'hd0bc; // 0x32e6
	13'h1974: q1 = 16'hffff; // 0x32e8
	13'h1975: q1 = 16'hffda; // 0x32ea
	13'h1976: q1 = 16'h2f00; // 0x32ec
	13'h1977: q1 = 16'h4eb9; // 0x32ee
	13'h1978: q1 = 16'h0000; // 0x32f0
	13'h1979: q1 = 16'h026c; // 0x32f2
	13'h197a: q1 = 16'hdefc; // 0x32f4
	13'h197b: q1 = 16'h000a; // 0x32f6
	13'h197c: q1 = 16'h4a79; // 0x32f8
	13'h197d: q1 = 16'h0001; // 0x32fa
	13'h197e: q1 = 16'h7582; // 0x32fc
	13'h197f: q1 = 16'h6f00; // 0x32fe
	13'h1980: q1 = 16'h00c0; // 0x3300
	13'h1981: q1 = 16'h3ebc; // 0x3302
	13'h1982: q1 = 16'h0013; // 0x3304
	13'h1983: q1 = 16'h200e; // 0x3306
	13'h1984: q1 = 16'hd0bc; // 0x3308
	13'h1985: q1 = 16'hffff; // 0x330a
	13'h1986: q1 = 16'hffda; // 0x330c
	13'h1987: q1 = 16'h2f00; // 0x330e
	13'h1988: q1 = 16'h4eb9; // 0x3310
	13'h1989: q1 = 16'h0000; // 0x3312
	13'h198a: q1 = 16'h78f6; // 0x3314
	13'h198b: q1 = 16'h4a9f; // 0x3316
	13'h198c: q1 = 16'h200e; // 0x3318
	13'h198d: q1 = 16'hd0bc; // 0x331a
	13'h198e: q1 = 16'hffff; // 0x331c
	13'h198f: q1 = 16'hffda; // 0x331e
	13'h1990: q1 = 16'h2e80; // 0x3320
	13'h1991: q1 = 16'h3f39; // 0x3322
	13'h1992: q1 = 16'h0001; // 0x3324
	13'h1993: q1 = 16'h7582; // 0x3326
	13'h1994: q1 = 16'h4eb9; // 0x3328
	13'h1995: q1 = 16'h0000; // 0x332a
	13'h1996: q1 = 16'h0798; // 0x332c
	13'h1997: q1 = 16'h4a5f; // 0x332e
	13'h1998: q1 = 16'h3ebc; // 0x3330
	13'h1999: q1 = 16'h0014; // 0x3332
	13'h199a: q1 = 16'h200e; // 0x3334
	13'h199b: q1 = 16'hd0bc; // 0x3336
	13'h199c: q1 = 16'hffff; // 0x3338
	13'h199d: q1 = 16'hffb8; // 0x333a
	13'h199e: q1 = 16'h2f00; // 0x333c
	13'h199f: q1 = 16'h4eb9; // 0x333e
	13'h19a0: q1 = 16'h0000; // 0x3340
	13'h19a1: q1 = 16'h78f6; // 0x3342
	13'h19a2: q1 = 16'h4a9f; // 0x3344
	13'h19a3: q1 = 16'h200e; // 0x3346
	13'h19a4: q1 = 16'hd0bc; // 0x3348
	13'h19a5: q1 = 16'hffff; // 0x334a
	13'h19a6: q1 = 16'hffb8; // 0x334c
	13'h19a7: q1 = 16'h2e80; // 0x334e
	13'h19a8: q1 = 16'h200e; // 0x3350
	13'h19a9: q1 = 16'hd0bc; // 0x3352
	13'h19aa: q1 = 16'hffff; // 0x3354
	13'h19ab: q1 = 16'hffda; // 0x3356
	13'h19ac: q1 = 16'h2f00; // 0x3358
	13'h19ad: q1 = 16'h4eb9; // 0x335a
	13'h19ae: q1 = 16'h0000; // 0x335c
	13'h19af: q1 = 16'h0770; // 0x335e
	13'h19b0: q1 = 16'h4a9f; // 0x3360
	13'h19b1: q1 = 16'h4a79; // 0x3362
	13'h19b2: q1 = 16'h0001; // 0x3364
	13'h19b3: q1 = 16'h7586; // 0x3366
	13'h19b4: q1 = 16'h6f32; // 0x3368
	13'h19b5: q1 = 16'h3ebc; // 0x336a
	13'h19b6: q1 = 16'h0015; // 0x336c
	13'h19b7: q1 = 16'h200e; // 0x336e
	13'h19b8: q1 = 16'hd0bc; // 0x3370
	13'h19b9: q1 = 16'hffff; // 0x3372
	13'h19ba: q1 = 16'hffb8; // 0x3374
	13'h19bb: q1 = 16'h2f00; // 0x3376
	13'h19bc: q1 = 16'h4eb9; // 0x3378
	13'h19bd: q1 = 16'h0000; // 0x337a
	13'h19be: q1 = 16'h78f6; // 0x337c
	13'h19bf: q1 = 16'h4a9f; // 0x337e
	13'h19c0: q1 = 16'h200e; // 0x3380
	13'h19c1: q1 = 16'hd0bc; // 0x3382
	13'h19c2: q1 = 16'hffff; // 0x3384
	13'h19c3: q1 = 16'hffb8; // 0x3386
	13'h19c4: q1 = 16'h2e80; // 0x3388
	13'h19c5: q1 = 16'h200e; // 0x338a
	13'h19c6: q1 = 16'hd0bc; // 0x338c
	13'h19c7: q1 = 16'hffff; // 0x338e
	13'h19c8: q1 = 16'hffda; // 0x3390
	13'h19c9: q1 = 16'h2f00; // 0x3392
	13'h19ca: q1 = 16'h4eb9; // 0x3394
	13'h19cb: q1 = 16'h0000; // 0x3396
	13'h19cc: q1 = 16'h0770; // 0x3398
	13'h19cd: q1 = 16'h4a9f; // 0x339a
	13'h19ce: q1 = 16'h3ebc; // 0x339c
	13'h19cf: q1 = 16'h002e; // 0x339e
	13'h19d0: q1 = 16'h3f3c; // 0x33a0
	13'h19d1: q1 = 16'h0020; // 0x33a2
	13'h19d2: q1 = 16'h3f3c; // 0x33a4
	13'h19d3: q1 = 16'h0064; // 0x33a6
	13'h19d4: q1 = 16'h3f06; // 0x33a8
	13'h19d5: q1 = 16'h5346; // 0x33aa
	13'h19d6: q1 = 16'h200e; // 0x33ac
	13'h19d7: q1 = 16'hd0bc; // 0x33ae
	13'h19d8: q1 = 16'hffff; // 0x33b0
	13'h19d9: q1 = 16'hffda; // 0x33b2
	13'h19da: q1 = 16'h2f00; // 0x33b4
	13'h19db: q1 = 16'h4eb9; // 0x33b6
	13'h19dc: q1 = 16'h0000; // 0x33b8
	13'h19dd: q1 = 16'h026c; // 0x33ba
	13'h19de: q1 = 16'hdefc; // 0x33bc
	13'h19df: q1 = 16'h000a; // 0x33be
	13'h19e0: q1 = 16'h4a79; // 0x33c0
	13'h19e1: q1 = 16'h0001; // 0x33c2
	13'h19e2: q1 = 16'h7586; // 0x33c4
	13'h19e3: q1 = 16'h6f6a; // 0x33c6
	13'h19e4: q1 = 16'h0c79; // 0x33c8
	13'h19e5: q1 = 16'h0003; // 0x33ca
	13'h19e6: q1 = 16'h0001; // 0x33cc
	13'h19e7: q1 = 16'h758c; // 0x33ce
	13'h19e8: q1 = 16'h6628; // 0x33d0
	13'h19e9: q1 = 16'h4a79; // 0x33d2
	13'h19ea: q1 = 16'h0001; // 0x33d4
	13'h19eb: q1 = 16'h7582; // 0x33d6
	13'h19ec: q1 = 16'h6620; // 0x33d8
	13'h19ed: q1 = 16'h3ebc; // 0x33da
	13'h19ee: q1 = 16'h002e; // 0x33dc
	13'h19ef: q1 = 16'h3f3c; // 0x33de
	13'h19f0: q1 = 16'h0020; // 0x33e0
	13'h19f1: q1 = 16'h3f3c; // 0x33e2
	13'h19f2: q1 = 16'h0064; // 0x33e4
	13'h19f3: q1 = 16'h3f06; // 0x33e6
	13'h19f4: q1 = 16'h5346; // 0x33e8
	13'h19f5: q1 = 16'h2f3c; // 0x33ea
	13'h19f6: q1 = 16'h0000; // 0x33ec
	13'h19f7: q1 = 16'hceb3; // 0x33ee
	13'h19f8: q1 = 16'h4eb9; // 0x33f0
	13'h19f9: q1 = 16'h0000; // 0x33f2
	13'h19fa: q1 = 16'h026c; // 0x33f4
	13'h19fb: q1 = 16'hdefc; // 0x33f6
	13'h19fc: q1 = 16'h000a; // 0x33f8
	13'h19fd: q1 = 16'h3ebc; // 0x33fa
	13'h19fe: q1 = 16'h0016; // 0x33fc
	13'h19ff: q1 = 16'h200e; // 0x33fe
	13'h1a00: q1 = 16'hd0bc; // 0x3400
	13'h1a01: q1 = 16'hffff; // 0x3402
	13'h1a02: q1 = 16'hffda; // 0x3404
	13'h1a03: q1 = 16'h2f00; // 0x3406
	13'h1a04: q1 = 16'h4eb9; // 0x3408
	13'h1a05: q1 = 16'h0000; // 0x340a
	13'h1a06: q1 = 16'h78f6; // 0x340c
	13'h1a07: q1 = 16'h4a9f; // 0x340e
	13'h1a08: q1 = 16'h3ebc; // 0x3410
	13'h1a09: q1 = 16'h0033; // 0x3412
	13'h1a0a: q1 = 16'h3f3c; // 0x3414
	13'h1a0b: q1 = 16'h0020; // 0x3416
	13'h1a0c: q1 = 16'h3f3c; // 0x3418
	13'h1a0d: q1 = 16'h0064; // 0x341a
	13'h1a0e: q1 = 16'h3f06; // 0x341c
	13'h1a0f: q1 = 16'h200e; // 0x341e
	13'h1a10: q1 = 16'hd0bc; // 0x3420
	13'h1a11: q1 = 16'hffff; // 0x3422
	13'h1a12: q1 = 16'hffda; // 0x3424
	13'h1a13: q1 = 16'h2f00; // 0x3426
	13'h1a14: q1 = 16'h4eb9; // 0x3428
	13'h1a15: q1 = 16'h0000; // 0x342a
	13'h1a16: q1 = 16'h026c; // 0x342c
	13'h1a17: q1 = 16'hdefc; // 0x342e
	13'h1a18: q1 = 16'h000a; // 0x3430
	13'h1a19: q1 = 16'h3ebc; // 0x3432
	13'h1a1a: q1 = 16'h0007; // 0x3434
	13'h1a1b: q1 = 16'h4eb9; // 0x3436
	13'h1a1c: q1 = 16'h0000; // 0x3438
	13'h1a1d: q1 = 16'h5be0; // 0x343a
	13'h1a1e: q1 = 16'h3ebc; // 0x343c
	13'h1a1f: q1 = 16'h0078; // 0x343e
	13'h1a20: q1 = 16'h4eb9; // 0x3440
	13'h1a21: q1 = 16'h0000; // 0x3442
	13'h1a22: q1 = 16'h6aca; // 0x3444
	13'h1a23: q1 = 16'h4a40; // 0x3446
	13'h1a24: q1 = 16'h33f9; // 0x3448
	13'h1a25: q1 = 16'h0001; // 0x344a
	13'h1a26: q1 = 16'h7eba; // 0x344c
	13'h1a27: q1 = 16'h0001; // 0x344e
	13'h1a28: q1 = 16'h8a76; // 0x3450
	13'h1a29: q1 = 16'h4279; // 0x3452
	13'h1a2a: q1 = 16'h0001; // 0x3454
	13'h1a2b: q1 = 16'h7faa; // 0x3456
	13'h1a2c: q1 = 16'h4279; // 0x3458
	13'h1a2d: q1 = 16'h0001; // 0x345a
	13'h1a2e: q1 = 16'h806e; // 0x345c
	13'h1a2f: q1 = 16'h4a9f; // 0x345e
	13'h1a30: q1 = 16'h4cdf; // 0x3460
	13'h1a31: q1 = 16'h30c0; // 0x3462
	13'h1a32: q1 = 16'h4e5e; // 0x3464
	13'h1a33: q1 = 16'h4e75; // 0x3466
	13'h1a34: q1 = 16'h4e56; // 0x3468
	13'h1a35: q1 = 16'hfffc; // 0x346a
	13'h1a36: q1 = 16'h48e7; // 0x346c
	13'h1a37: q1 = 16'h0304; // 0x346e
	13'h1a38: q1 = 16'h4ab9; // 0x3470
	13'h1a39: q1 = 16'h0001; // 0x3472
	13'h1a3a: q1 = 16'h7fa2; // 0x3474
	13'h1a3b: q1 = 16'h6f06; // 0x3476
	13'h1a3c: q1 = 16'h53b9; // 0x3478
	13'h1a3d: q1 = 16'h0001; // 0x347a
	13'h1a3e: q1 = 16'h7fa2; // 0x347c
	13'h1a3f: q1 = 16'h4ab9; // 0x347e
	13'h1a40: q1 = 16'h0001; // 0x3480
	13'h1a41: q1 = 16'h7f60; // 0x3482
	13'h1a42: q1 = 16'h6f06; // 0x3484
	13'h1a43: q1 = 16'h53b9; // 0x3486
	13'h1a44: q1 = 16'h0001; // 0x3488
	13'h1a45: q1 = 16'h7f60; // 0x348a
	13'h1a46: q1 = 16'h4ab9; // 0x348c
	13'h1a47: q1 = 16'h0001; // 0x348e
	13'h1a48: q1 = 16'h7fc2; // 0x3490
	13'h1a49: q1 = 16'h6f06; // 0x3492
	13'h1a4a: q1 = 16'h53b9; // 0x3494
	13'h1a4b: q1 = 16'h0001; // 0x3496
	13'h1a4c: q1 = 16'h7fc2; // 0x3498
	13'h1a4d: q1 = 16'h4ab9; // 0x349a
	13'h1a4e: q1 = 16'h0001; // 0x349c
	13'h1a4f: q1 = 16'h7fac; // 0x349e
	13'h1a50: q1 = 16'h6f06; // 0x34a0
	13'h1a51: q1 = 16'h53b9; // 0x34a2
	13'h1a52: q1 = 16'h0001; // 0x34a4
	13'h1a53: q1 = 16'h7fac; // 0x34a6
	13'h1a54: q1 = 16'h4a79; // 0x34a8
	13'h1a55: q1 = 16'h0001; // 0x34aa
	13'h1a56: q1 = 16'h7fb0; // 0x34ac
	13'h1a57: q1 = 16'h6f08; // 0x34ae
	13'h1a58: q1 = 16'h5379; // 0x34b0
	13'h1a59: q1 = 16'h0001; // 0x34b2
	13'h1a5a: q1 = 16'h7fb0; // 0x34b4
	13'h1a5b: q1 = 16'h6014; // 0x34b6
	13'h1a5c: q1 = 16'h33fc; // 0x34b8
	13'h1a5d: q1 = 16'h003c; // 0x34ba
	13'h1a5e: q1 = 16'h0001; // 0x34bc
	13'h1a5f: q1 = 16'h7fb0; // 0x34be
	13'h1a60: q1 = 16'h52b9; // 0x34c0
	13'h1a61: q1 = 16'h0001; // 0x34c2
	13'h1a62: q1 = 16'h75d2; // 0x34c4
	13'h1a63: q1 = 16'h52b9; // 0x34c6
	13'h1a64: q1 = 16'h0001; // 0x34c8
	13'h1a65: q1 = 16'h75ca; // 0x34ca
	13'h1a66: q1 = 16'h52b9; // 0x34cc
	13'h1a67: q1 = 16'h0001; // 0x34ce
	13'h1a68: q1 = 16'h7596; // 0x34d0
	13'h1a69: q1 = 16'h2a79; // 0x34d2
	13'h1a6a: q1 = 16'h0000; // 0x34d4
	13'h1a6b: q1 = 16'hceb8; // 0x34d6
	13'h1a6c: q1 = 16'h3e15; // 0x34d8
	13'h1a6d: q1 = 16'h2a79; // 0x34da
	13'h1a6e: q1 = 16'h0000; // 0x34dc
	13'h1a6f: q1 = 16'hcebc; // 0x34de
	13'h1a70: q1 = 16'h3e15; // 0x34e0
	13'h1a71: q1 = 16'h4a79; // 0x34e2
	13'h1a72: q1 = 16'h0001; // 0x34e4
	13'h1a73: q1 = 16'h8052; // 0x34e6
	13'h1a74: q1 = 16'h6714; // 0x34e8
	13'h1a75: q1 = 16'h0807; // 0x34ea
	13'h1a76: q1 = 16'h0006; // 0x34ec
	13'h1a77: q1 = 16'h6704; // 0x34ee
	13'h1a78: q1 = 16'h4240; // 0x34f0
	13'h1a79: q1 = 16'h6002; // 0x34f2
	13'h1a7a: q1 = 16'h7001; // 0x34f4
	13'h1a7b: q1 = 16'h33c0; // 0x34f6
	13'h1a7c: q1 = 16'h0001; // 0x34f8
	13'h1a7d: q1 = 16'h7fca; // 0x34fa
	13'h1a7e: q1 = 16'h6012; // 0x34fc
	13'h1a7f: q1 = 16'h0807; // 0x34fe
	13'h1a80: q1 = 16'h0005; // 0x3500
	13'h1a81: q1 = 16'h6704; // 0x3502
	13'h1a82: q1 = 16'h4240; // 0x3504
	13'h1a83: q1 = 16'h6002; // 0x3506
	13'h1a84: q1 = 16'h7001; // 0x3508
	13'h1a85: q1 = 16'h33c0; // 0x350a
	13'h1a86: q1 = 16'h0001; // 0x350c
	13'h1a87: q1 = 16'h7fca; // 0x350e
	13'h1a88: q1 = 16'h0807; // 0x3510
	13'h1a89: q1 = 16'h0002; // 0x3512
	13'h1a8a: q1 = 16'h6704; // 0x3514
	13'h1a8b: q1 = 16'h4240; // 0x3516
	13'h1a8c: q1 = 16'h6002; // 0x3518
	13'h1a8d: q1 = 16'h7001; // 0x351a
	13'h1a8e: q1 = 16'h33c0; // 0x351c
	13'h1a8f: q1 = 16'h0001; // 0x351e
	13'h1a90: q1 = 16'h8a7e; // 0x3520
	13'h1a91: q1 = 16'h0807; // 0x3522
	13'h1a92: q1 = 16'h0003; // 0x3524
	13'h1a93: q1 = 16'h6704; // 0x3526
	13'h1a94: q1 = 16'h4240; // 0x3528
	13'h1a95: q1 = 16'h6002; // 0x352a
	13'h1a96: q1 = 16'h7001; // 0x352c
	13'h1a97: q1 = 16'h33c0; // 0x352e
	13'h1a98: q1 = 16'h0001; // 0x3530
	13'h1a99: q1 = 16'h8a80; // 0x3532
	13'h1a9a: q1 = 16'h4279; // 0x3534
	13'h1a9b: q1 = 16'h0001; // 0x3536
	13'h1a9c: q1 = 16'h7f5e; // 0x3538
	13'h1a9d: q1 = 16'h4a79; // 0x353a
	13'h1a9e: q1 = 16'h0001; // 0x353c
	13'h1a9f: q1 = 16'h8a7e; // 0x353e
	13'h1aa0: q1 = 16'h6712; // 0x3540
	13'h1aa1: q1 = 16'h4a79; // 0x3542
	13'h1aa2: q1 = 16'h0001; // 0x3544
	13'h1aa3: q1 = 16'h7594; // 0x3546
	13'h1aa4: q1 = 16'h670a; // 0x3548
	13'h1aa5: q1 = 16'h33fc; // 0x354a
	13'h1aa6: q1 = 16'h0001; // 0x354c
	13'h1aa7: q1 = 16'h0001; // 0x354e
	13'h1aa8: q1 = 16'h7f5e; // 0x3550
	13'h1aa9: q1 = 16'h601a; // 0x3552
	13'h1aaa: q1 = 16'h4a79; // 0x3554
	13'h1aab: q1 = 16'h0001; // 0x3556
	13'h1aac: q1 = 16'h8a80; // 0x3558
	13'h1aad: q1 = 16'h6712; // 0x355a
	13'h1aae: q1 = 16'h0c79; // 0x355c
	13'h1aaf: q1 = 16'h0001; // 0x355e
	13'h1ab0: q1 = 16'h0001; // 0x3560
	13'h1ab1: q1 = 16'h7594; // 0x3562
	13'h1ab2: q1 = 16'h6f08; // 0x3564
	13'h1ab3: q1 = 16'h33fc; // 0x3566
	13'h1ab4: q1 = 16'h0002; // 0x3568
	13'h1ab5: q1 = 16'h0001; // 0x356a
	13'h1ab6: q1 = 16'h7f5e; // 0x356c
	13'h1ab7: q1 = 16'h0807; // 0x356e
	13'h1ab8: q1 = 16'h0007; // 0x3570
	13'h1ab9: q1 = 16'h6704; // 0x3572
	13'h1aba: q1 = 16'h4240; // 0x3574
	13'h1abb: q1 = 16'h6002; // 0x3576
	13'h1abc: q1 = 16'h7001; // 0x3578
	13'h1abd: q1 = 16'h33c0; // 0x357a
	13'h1abe: q1 = 16'h0001; // 0x357c
	13'h1abf: q1 = 16'h8a7c; // 0x357e
	13'h1ac0: q1 = 16'h2a79; // 0x3580
	13'h1ac1: q1 = 16'h0000; // 0x3582
	13'h1ac2: q1 = 16'hcec0; // 0x3584
	13'h1ac3: q1 = 16'h302d; // 0x3586
	13'h1ac4: q1 = 16'h0010; // 0x3588
	13'h1ac5: q1 = 16'hc07c; // 0x358a
	13'h1ac6: q1 = 16'h00ff; // 0x358c
	13'h1ac7: q1 = 16'h663c; // 0x358e
	13'h1ac8: q1 = 16'h4247; // 0x3590
	13'h1ac9: q1 = 16'hbe7c; // 0x3592
	13'h1aca: q1 = 16'h0008; // 0x3594
	13'h1acb: q1 = 16'h6c28; // 0x3596
	13'h1acc: q1 = 16'h7007; // 0x3598
	13'h1acd: q1 = 16'h9047; // 0x359a
	13'h1ace: q1 = 16'he340; // 0x359c
	13'h1acf: q1 = 16'h48c0; // 0x359e
	13'h1ad0: q1 = 16'hd0bc; // 0x35a0
	13'h1ad1: q1 = 16'h0001; // 0x35a2
	13'h1ad2: q1 = 16'h805c; // 0x35a4
	13'h1ad3: q1 = 16'h2040; // 0x35a6
	13'h1ad4: q1 = 16'h3207; // 0x35a8
	13'h1ad5: q1 = 16'he341; // 0x35aa
	13'h1ad6: q1 = 16'h48c1; // 0x35ac
	13'h1ad7: q1 = 16'hd28d; // 0x35ae
	13'h1ad8: q1 = 16'h2241; // 0x35b0
	13'h1ad9: q1 = 16'h3211; // 0x35b2
	13'h1ada: q1 = 16'hc27c; // 0x35b4
	13'h1adb: q1 = 16'h00ff; // 0x35b6
	13'h1adc: q1 = 16'hee41; // 0x35b8
	13'h1add: q1 = 16'h3081; // 0x35ba
	13'h1ade: q1 = 16'h5247; // 0x35bc
	13'h1adf: q1 = 16'h60d2; // 0x35be
	13'h1ae0: q1 = 16'h3b7c; // 0x35c0
	13'h1ae1: q1 = 16'h0003; // 0x35c2
	13'h1ae2: q1 = 16'h001e; // 0x35c4
	13'h1ae3: q1 = 16'h3b7c; // 0x35c6
	13'h1ae4: q1 = 16'h0007; // 0x35c8
	13'h1ae5: q1 = 16'h0016; // 0x35ca
	13'h1ae6: q1 = 16'h3e39; // 0x35cc
	13'h1ae7: q1 = 16'h0001; // 0x35ce
	13'h1ae8: q1 = 16'h861e; // 0x35d0
	13'h1ae9: q1 = 16'h4a79; // 0x35d2
	13'h1aea: q1 = 16'h0001; // 0x35d4
	13'h1aeb: q1 = 16'h8a7c; // 0x35d6
	13'h1aec: q1 = 16'h6626; // 0x35d8
	13'h1aed: q1 = 16'h4a79; // 0x35da
	13'h1aee: q1 = 16'h0001; // 0x35dc
	13'h1aef: q1 = 16'h867a; // 0x35de
	13'h1af0: q1 = 16'h671e; // 0x35e0
	13'h1af1: q1 = 16'h0c79; // 0x35e2
	13'h1af2: q1 = 16'h0001; // 0x35e4
	13'h1af3: q1 = 16'h0001; // 0x35e6
	13'h1af4: q1 = 16'h87dc; // 0x35e8
	13'h1af5: q1 = 16'h660a; // 0x35ea
	13'h1af6: q1 = 16'hce7c; // 0x35ec
	13'h1af7: q1 = 16'hffdf; // 0x35ee
	13'h1af8: q1 = 16'h8e7c; // 0x35f0
	13'h1af9: q1 = 16'h0010; // 0x35f2
	13'h1afa: q1 = 16'h6008; // 0x35f4
	13'h1afb: q1 = 16'hce7c; // 0x35f6
	13'h1afc: q1 = 16'hffef; // 0x35f8
	13'h1afd: q1 = 16'h8e7c; // 0x35fa
	13'h1afe: q1 = 16'h0020; // 0x35fc
	13'h1aff: q1 = 16'h6032; // 0x35fe
	13'h1b00: q1 = 16'h4a79; // 0x3600
	13'h1b01: q1 = 16'h0001; // 0x3602
	13'h1b02: q1 = 16'h8a7c; // 0x3604
	13'h1b03: q1 = 16'h6626; // 0x3606
	13'h1b04: q1 = 16'h4a79; // 0x3608
	13'h1b05: q1 = 16'h0001; // 0x360a
	13'h1b06: q1 = 16'h7594; // 0x360c
	13'h1b07: q1 = 16'h671e; // 0x360e
	13'h1b08: q1 = 16'h0c79; // 0x3610
	13'h1b09: q1 = 16'h001e; // 0x3612
	13'h1b0a: q1 = 16'h0001; // 0x3614
	13'h1b0b: q1 = 16'h7fb0; // 0x3616
	13'h1b0c: q1 = 16'h6c14; // 0x3618
	13'h1b0d: q1 = 16'h8e7c; // 0x361a
	13'h1b0e: q1 = 16'h0010; // 0x361c
	13'h1b0f: q1 = 16'h0c79; // 0x361e
	13'h1b10: q1 = 16'h0001; // 0x3620
	13'h1b11: q1 = 16'h0001; // 0x3622
	13'h1b12: q1 = 16'h7594; // 0x3624
	13'h1b13: q1 = 16'h6f04; // 0x3626
	13'h1b14: q1 = 16'h8e7c; // 0x3628
	13'h1b15: q1 = 16'h0020; // 0x362a
	13'h1b16: q1 = 16'h6004; // 0x362c
	13'h1b17: q1 = 16'hce7c; // 0x362e
	13'h1b18: q1 = 16'hffcf; // 0x3630
	13'h1b19: q1 = 16'h4a79; // 0x3632
	13'h1b1a: q1 = 16'h0001; // 0x3634
	13'h1b1b: q1 = 16'h7fa6; // 0x3636
	13'h1b1c: q1 = 16'h6706; // 0x3638
	13'h1b1d: q1 = 16'h8e7c; // 0x363a
	13'h1b1e: q1 = 16'h0001; // 0x363c
	13'h1b1f: q1 = 16'h6004; // 0x363e
	13'h1b20: q1 = 16'hce7c; // 0x3640
	13'h1b21: q1 = 16'hfffe; // 0x3642
	13'h1b22: q1 = 16'hce7c; // 0x3644
	13'h1b23: q1 = 16'hff3f; // 0x3646
	13'h1b24: q1 = 16'h4a79; // 0x3648
	13'h1b25: q1 = 16'h0001; // 0x364a
	13'h1b26: q1 = 16'h867c; // 0x364c
	13'h1b27: q1 = 16'h6706; // 0x364e
	13'h1b28: q1 = 16'h303c; // 0x3650
	13'h1b29: q1 = 16'h0080; // 0x3652
	13'h1b2a: q1 = 16'h6002; // 0x3654
	13'h1b2b: q1 = 16'h4240; // 0x3656
	13'h1b2c: q1 = 16'h4a79; // 0x3658
	13'h1b2d: q1 = 16'h0001; // 0x365a
	13'h1b2e: q1 = 16'h861a; // 0x365c
	13'h1b2f: q1 = 16'h6704; // 0x365e
	13'h1b30: q1 = 16'h7240; // 0x3660
	13'h1b31: q1 = 16'h6002; // 0x3662
	13'h1b32: q1 = 16'h4241; // 0x3664
	13'h1b33: q1 = 16'h8041; // 0x3666
	13'h1b34: q1 = 16'h8e40; // 0x3668
	13'h1b35: q1 = 16'h4a79; // 0x366a
	13'h1b36: q1 = 16'h0001; // 0x366c
	13'h1b37: q1 = 16'h867c; // 0x366e
	13'h1b38: q1 = 16'h6706; // 0x3670
	13'h1b39: q1 = 16'h5379; // 0x3672
	13'h1b3a: q1 = 16'h0001; // 0x3674
	13'h1b3b: q1 = 16'h867c; // 0x3676
	13'h1b3c: q1 = 16'h4a79; // 0x3678
	13'h1b3d: q1 = 16'h0001; // 0x367a
	13'h1b3e: q1 = 16'h861a; // 0x367c
	13'h1b3f: q1 = 16'h6706; // 0x367e
	13'h1b40: q1 = 16'h5379; // 0x3680
	13'h1b41: q1 = 16'h0001; // 0x3682
	13'h1b42: q1 = 16'h861a; // 0x3684
	13'h1b43: q1 = 16'h33c7; // 0x3686
	13'h1b44: q1 = 16'h0001; // 0x3688
	13'h1b45: q1 = 16'h861e; // 0x368a
	13'h1b46: q1 = 16'h2a79; // 0x368c
	13'h1b47: q1 = 16'h0000; // 0x368e
	13'h1b48: q1 = 16'hcebc; // 0x3690
	13'h1b49: q1 = 16'h3ab9; // 0x3692
	13'h1b4a: q1 = 16'h0001; // 0x3694
	13'h1b4b: q1 = 16'h861e; // 0x3696
	13'h1b4c: q1 = 16'h2a79; // 0x3698
	13'h1b4d: q1 = 16'h0000; // 0x369a
	13'h1b4e: q1 = 16'hcec4; // 0x369c
	13'h1b4f: q1 = 16'h3e15; // 0x369e
	13'h1b50: q1 = 16'h4a79; // 0x36a0
	13'h1b51: q1 = 16'h0001; // 0x36a2
	13'h1b52: q1 = 16'h7fcc; // 0x36a4
	13'h1b53: q1 = 16'h670e; // 0x36a6
	13'h1b54: q1 = 16'h3007; // 0x36a8
	13'h1b55: q1 = 16'hc07c; // 0x36aa
	13'h1b56: q1 = 16'h00ff; // 0x36ac
	13'h1b57: q1 = 16'h33c0; // 0x36ae
	13'h1b58: q1 = 16'h0001; // 0x36b0
	13'h1b59: q1 = 16'h861c; // 0x36b2
	13'h1b5a: q1 = 16'h600c; // 0x36b4
	13'h1b5b: q1 = 16'h3007; // 0x36b6
	13'h1b5c: q1 = 16'hc07c; // 0x36b8
	13'h1b5d: q1 = 16'h00ff; // 0x36ba
	13'h1b5e: q1 = 16'h33c0; // 0x36bc
	13'h1b5f: q1 = 16'h0001; // 0x36be
	13'h1b60: q1 = 16'h8626; // 0x36c0
	13'h1b61: q1 = 16'h4a79; // 0x36c2
	13'h1b62: q1 = 16'h0001; // 0x36c4
	13'h1b63: q1 = 16'h7fcc; // 0x36c6
	13'h1b64: q1 = 16'h6714; // 0x36c8
	13'h1b65: q1 = 16'h4a79; // 0x36ca
	13'h1b66: q1 = 16'h0001; // 0x36cc
	13'h1b67: q1 = 16'h7fbe; // 0x36ce
	13'h1b68: q1 = 16'h670c; // 0x36d0
	13'h1b69: q1 = 16'h33f9; // 0x36d2
	13'h1b6a: q1 = 16'h0001; // 0x36d4
	13'h1b6b: q1 = 16'h861c; // 0x36d6
	13'h1b6c: q1 = 16'h0001; // 0x36d8
	13'h1b6d: q1 = 16'h86b4; // 0x36da
	13'h1b6e: q1 = 16'h6042; // 0x36dc
	13'h1b6f: q1 = 16'h4a79; // 0x36de
	13'h1b70: q1 = 16'h0001; // 0x36e0
	13'h1b71: q1 = 16'h7fcc; // 0x36e2
	13'h1b72: q1 = 16'h6714; // 0x36e4
	13'h1b73: q1 = 16'h4a79; // 0x36e6
	13'h1b74: q1 = 16'h0001; // 0x36e8
	13'h1b75: q1 = 16'h7fbe; // 0x36ea
	13'h1b76: q1 = 16'h660c; // 0x36ec
	13'h1b77: q1 = 16'h33f9; // 0x36ee
	13'h1b78: q1 = 16'h0001; // 0x36f0
	13'h1b79: q1 = 16'h861c; // 0x36f2
	13'h1b7a: q1 = 16'h0001; // 0x36f4
	13'h1b7b: q1 = 16'h86b2; // 0x36f6
	13'h1b7c: q1 = 16'h6026; // 0x36f8
	13'h1b7d: q1 = 16'h4a79; // 0x36fa
	13'h1b7e: q1 = 16'h0001; // 0x36fc
	13'h1b7f: q1 = 16'h7fcc; // 0x36fe
	13'h1b80: q1 = 16'h6614; // 0x3700
	13'h1b81: q1 = 16'h4a79; // 0x3702
	13'h1b82: q1 = 16'h0001; // 0x3704
	13'h1b83: q1 = 16'h7fbe; // 0x3706
	13'h1b84: q1 = 16'h670c; // 0x3708
	13'h1b85: q1 = 16'h33f9; // 0x370a
	13'h1b86: q1 = 16'h0001; // 0x370c
	13'h1b87: q1 = 16'h8626; // 0x370e
	13'h1b88: q1 = 16'h0001; // 0x3710
	13'h1b89: q1 = 16'h86da; // 0x3712
	13'h1b8a: q1 = 16'h600a; // 0x3714
	13'h1b8b: q1 = 16'h33f9; // 0x3716
	13'h1b8c: q1 = 16'h0001; // 0x3718
	13'h1b8d: q1 = 16'h8626; // 0x371a
	13'h1b8e: q1 = 16'h0001; // 0x371c
	13'h1b8f: q1 = 16'h86b6; // 0x371e
	13'h1b90: q1 = 16'h4a79; // 0x3720
	13'h1b91: q1 = 16'h0001; // 0x3722
	13'h1b92: q1 = 16'h8052; // 0x3724
	13'h1b93: q1 = 16'h6720; // 0x3726
	13'h1b94: q1 = 16'h4a79; // 0x3728
	13'h1b95: q1 = 16'h0001; // 0x372a
	13'h1b96: q1 = 16'h7fcc; // 0x372c
	13'h1b97: q1 = 16'h6708; // 0x372e
	13'h1b98: q1 = 16'h2a79; // 0x3730
	13'h1b99: q1 = 16'h0000; // 0x3732
	13'h1b9a: q1 = 16'hcec8; // 0x3734
	13'h1b9b: q1 = 16'h6006; // 0x3736
	13'h1b9c: q1 = 16'h2a79; // 0x3738
	13'h1b9d: q1 = 16'h0000; // 0x373a
	13'h1b9e: q1 = 16'hcecc; // 0x373c
	13'h1b9f: q1 = 16'h33fc; // 0x373e
	13'h1ba0: q1 = 16'h0001; // 0x3740
	13'h1ba1: q1 = 16'h0001; // 0x3742
	13'h1ba2: q1 = 16'h7fbe; // 0x3744
	13'h1ba3: q1 = 16'h601c; // 0x3746
	13'h1ba4: q1 = 16'h4a79; // 0x3748
	13'h1ba5: q1 = 16'h0001; // 0x374a
	13'h1ba6: q1 = 16'h7fcc; // 0x374c
	13'h1ba7: q1 = 16'h6708; // 0x374e
	13'h1ba8: q1 = 16'h2a79; // 0x3750
	13'h1ba9: q1 = 16'h0000; // 0x3752
	13'h1baa: q1 = 16'hced0; // 0x3754
	13'h1bab: q1 = 16'h6006; // 0x3756
	13'h1bac: q1 = 16'h2a79; // 0x3758
	13'h1bad: q1 = 16'h0000; // 0x375a
	13'h1bae: q1 = 16'hced4; // 0x375c
	13'h1baf: q1 = 16'h4279; // 0x375e
	13'h1bb0: q1 = 16'h0001; // 0x3760
	13'h1bb1: q1 = 16'h7fbe; // 0x3762
	13'h1bb2: q1 = 16'h3a87; // 0x3764
	13'h1bb3: q1 = 16'h2a79; // 0x3766
	13'h1bb4: q1 = 16'h0000; // 0x3768
	13'h1bb5: q1 = 16'hced8; // 0x376a
	13'h1bb6: q1 = 16'h3e15; // 0x376c
	13'h1bb7: q1 = 16'h7001; // 0x376e
	13'h1bb8: q1 = 16'h9079; // 0x3770
	13'h1bb9: q1 = 16'h0001; // 0x3772
	13'h1bba: q1 = 16'h7fcc; // 0x3774
	13'h1bbb: q1 = 16'h33c0; // 0x3776
	13'h1bbc: q1 = 16'h0001; // 0x3778
	13'h1bbd: q1 = 16'h7fcc; // 0x377a
	13'h1bbe: q1 = 16'h3039; // 0x377c
	13'h1bbf: q1 = 16'h0001; // 0x377e
	13'h1bc0: q1 = 16'h8052; // 0x3780
	13'h1bc1: q1 = 16'he740; // 0x3782
	13'h1bc2: q1 = 16'h48c0; // 0x3784
	13'h1bc3: q1 = 16'hd0bc; // 0x3786
	13'h1bc4: q1 = 16'h0001; // 0x3788
	13'h1bc5: q1 = 16'h8684; // 0x378a
	13'h1bc6: q1 = 16'h23c0; // 0x378c
	13'h1bc7: q1 = 16'h0001; // 0x378e
	13'h1bc8: q1 = 16'h7eb2; // 0x3790
	13'h1bc9: q1 = 16'h4a79; // 0x3792
	13'h1bca: q1 = 16'h0001; // 0x3794
	13'h1bcb: q1 = 16'h7fcc; // 0x3796
	13'h1bcc: q1 = 16'h6600; // 0x3798
	13'h1bcd: q1 = 16'h0078; // 0x379a
	13'h1bce: q1 = 16'h3039; // 0x379c
	13'h1bcf: q1 = 16'h0001; // 0x379e
	13'h1bd0: q1 = 16'h861c; // 0x37a0
	13'h1bd1: q1 = 16'hb079; // 0x37a2
	13'h1bd2: q1 = 16'h0001; // 0x37a4
	13'h1bd3: q1 = 16'h86d8; // 0x37a6
	13'h1bd4: q1 = 16'h6654; // 0x37a8
	13'h1bd5: q1 = 16'h5279; // 0x37aa
	13'h1bd6: q1 = 16'h0001; // 0x37ac
	13'h1bd7: q1 = 16'h8680; // 0x37ae
	13'h1bd8: q1 = 16'h0c79; // 0x37b0
	13'h1bd9: q1 = 16'h0005; // 0x37b2
	13'h1bda: q1 = 16'h0001; // 0x37b4
	13'h1bdb: q1 = 16'h8680; // 0x37b6
	13'h1bdc: q1 = 16'h6642; // 0x37b8
	13'h1bdd: q1 = 16'h2079; // 0x37ba
	13'h1bde: q1 = 16'h0001; // 0x37bc
	13'h1bdf: q1 = 16'h7eb2; // 0x37be
	13'h1be0: q1 = 16'h3010; // 0x37c0
	13'h1be1: q1 = 16'hb079; // 0x37c2
	13'h1be2: q1 = 16'h0001; // 0x37c4
	13'h1be3: q1 = 16'h861c; // 0x37c6
	13'h1be4: q1 = 16'h6f0c; // 0x37c8
	13'h1be5: q1 = 16'h2079; // 0x37ca
	13'h1be6: q1 = 16'h0001; // 0x37cc
	13'h1be7: q1 = 16'h7eb2; // 0x37ce
	13'h1be8: q1 = 16'h30b9; // 0x37d0
	13'h1be9: q1 = 16'h0001; // 0x37d2
	13'h1bea: q1 = 16'h861c; // 0x37d4
	13'h1beb: q1 = 16'h2079; // 0x37d6
	13'h1bec: q1 = 16'h0001; // 0x37d8
	13'h1bed: q1 = 16'h7eb2; // 0x37da
	13'h1bee: q1 = 16'h3028; // 0x37dc
	13'h1bef: q1 = 16'h0002; // 0x37de
	13'h1bf0: q1 = 16'hb079; // 0x37e0
	13'h1bf1: q1 = 16'h0001; // 0x37e2
	13'h1bf2: q1 = 16'h861c; // 0x37e4
	13'h1bf3: q1 = 16'h6c0e; // 0x37e6
	13'h1bf4: q1 = 16'h2079; // 0x37e8
	13'h1bf5: q1 = 16'h0001; // 0x37ea
	13'h1bf6: q1 = 16'h7eb2; // 0x37ec
	13'h1bf7: q1 = 16'h3179; // 0x37ee
	13'h1bf8: q1 = 16'h0001; // 0x37f0
	13'h1bf9: q1 = 16'h861c; // 0x37f2
	13'h1bfa: q1 = 16'h0002; // 0x37f4
	13'h1bfb: q1 = 16'h4279; // 0x37f6
	13'h1bfc: q1 = 16'h0001; // 0x37f8
	13'h1bfd: q1 = 16'h8680; // 0x37fa
	13'h1bfe: q1 = 16'h6006; // 0x37fc
	13'h1bff: q1 = 16'h4279; // 0x37fe
	13'h1c00: q1 = 16'h0001; // 0x3800
	13'h1c01: q1 = 16'h8680; // 0x3802
	13'h1c02: q1 = 16'h33f9; // 0x3804
	13'h1c03: q1 = 16'h0001; // 0x3806
	13'h1c04: q1 = 16'h861c; // 0x3808
	13'h1c05: q1 = 16'h0001; // 0x380a
	13'h1c06: q1 = 16'h86d8; // 0x380c
	13'h1c07: q1 = 16'h6000; // 0x380e
	13'h1c08: q1 = 16'h0078; // 0x3810
	13'h1c09: q1 = 16'h3039; // 0x3812
	13'h1c0a: q1 = 16'h0001; // 0x3814
	13'h1c0b: q1 = 16'h8626; // 0x3816
	13'h1c0c: q1 = 16'hb079; // 0x3818
	13'h1c0d: q1 = 16'h0001; // 0x381a
	13'h1c0e: q1 = 16'h87de; // 0x381c
	13'h1c0f: q1 = 16'h6658; // 0x381e
	13'h1c10: q1 = 16'h5279; // 0x3820
	13'h1c11: q1 = 16'h0001; // 0x3822
	13'h1c12: q1 = 16'h86aa; // 0x3824
	13'h1c13: q1 = 16'h0c79; // 0x3826
	13'h1c14: q1 = 16'h0005; // 0x3828
	13'h1c15: q1 = 16'h0001; // 0x382a
	13'h1c16: q1 = 16'h86aa; // 0x382c
	13'h1c17: q1 = 16'h6646; // 0x382e
	13'h1c18: q1 = 16'h2079; // 0x3830
	13'h1c19: q1 = 16'h0001; // 0x3832
	13'h1c1a: q1 = 16'h7eb2; // 0x3834
	13'h1c1b: q1 = 16'h3028; // 0x3836
	13'h1c1c: q1 = 16'h0004; // 0x3838
	13'h1c1d: q1 = 16'hb079; // 0x383a
	13'h1c1e: q1 = 16'h0001; // 0x383c
	13'h1c1f: q1 = 16'h8626; // 0x383e
	13'h1c20: q1 = 16'h6f0e; // 0x3840
	13'h1c21: q1 = 16'h2079; // 0x3842
	13'h1c22: q1 = 16'h0001; // 0x3844
	13'h1c23: q1 = 16'h7eb2; // 0x3846
	13'h1c24: q1 = 16'h3179; // 0x3848
	13'h1c25: q1 = 16'h0001; // 0x384a
	13'h1c26: q1 = 16'h8626; // 0x384c
	13'h1c27: q1 = 16'h0004; // 0x384e
	13'h1c28: q1 = 16'h2079; // 0x3850
	13'h1c29: q1 = 16'h0001; // 0x3852
	13'h1c2a: q1 = 16'h7eb2; // 0x3854
	13'h1c2b: q1 = 16'h3028; // 0x3856
	13'h1c2c: q1 = 16'h0006; // 0x3858
	13'h1c2d: q1 = 16'hb079; // 0x385a
	13'h1c2e: q1 = 16'h0001; // 0x385c
	13'h1c2f: q1 = 16'h8626; // 0x385e
	13'h1c30: q1 = 16'h6c0e; // 0x3860
	13'h1c31: q1 = 16'h2079; // 0x3862
	13'h1c32: q1 = 16'h0001; // 0x3864
	13'h1c33: q1 = 16'h7eb2; // 0x3866
	13'h1c34: q1 = 16'h3179; // 0x3868
	13'h1c35: q1 = 16'h0001; // 0x386a
	13'h1c36: q1 = 16'h8626; // 0x386c
	13'h1c37: q1 = 16'h0006; // 0x386e
	13'h1c38: q1 = 16'h4279; // 0x3870
	13'h1c39: q1 = 16'h0001; // 0x3872
	13'h1c3a: q1 = 16'h86aa; // 0x3874
	13'h1c3b: q1 = 16'h6006; // 0x3876
	13'h1c3c: q1 = 16'h4279; // 0x3878
	13'h1c3d: q1 = 16'h0001; // 0x387a
	13'h1c3e: q1 = 16'h86aa; // 0x387c
	13'h1c3f: q1 = 16'h33f9; // 0x387e
	13'h1c40: q1 = 16'h0001; // 0x3880
	13'h1c41: q1 = 16'h8626; // 0x3882
	13'h1c42: q1 = 16'h0001; // 0x3884
	13'h1c43: q1 = 16'h87de; // 0x3886
	13'h1c44: q1 = 16'h2079; // 0x3888
	13'h1c45: q1 = 16'h0001; // 0x388a
	13'h1c46: q1 = 16'h7eb2; // 0x388c
	13'h1c47: q1 = 16'h3028; // 0x388e
	13'h1c48: q1 = 16'h0002; // 0x3890
	13'h1c49: q1 = 16'h2279; // 0x3892
	13'h1c4a: q1 = 16'h0001; // 0x3894
	13'h1c4b: q1 = 16'h7eb2; // 0x3896
	13'h1c4c: q1 = 16'h9051; // 0x3898
	13'h1c4d: q1 = 16'he240; // 0x389a
	13'h1c4e: q1 = 16'h2279; // 0x389c
	13'h1c4f: q1 = 16'h0001; // 0x389e
	13'h1c50: q1 = 16'h7eb2; // 0x38a0
	13'h1c51: q1 = 16'hd051; // 0x38a2
	13'h1c52: q1 = 16'h3d40; // 0x38a4
	13'h1c53: q1 = 16'hfffe; // 0x38a6
	13'h1c54: q1 = 16'h2079; // 0x38a8
	13'h1c55: q1 = 16'h0001; // 0x38aa
	13'h1c56: q1 = 16'h7eb2; // 0x38ac
	13'h1c57: q1 = 16'h3028; // 0x38ae
	13'h1c58: q1 = 16'h0006; // 0x38b0
	13'h1c59: q1 = 16'h2279; // 0x38b2
	13'h1c5a: q1 = 16'h0001; // 0x38b4
	13'h1c5b: q1 = 16'h7eb2; // 0x38b6
	13'h1c5c: q1 = 16'h9069; // 0x38b8
	13'h1c5d: q1 = 16'h0004; // 0x38ba
	13'h1c5e: q1 = 16'he240; // 0x38bc
	13'h1c5f: q1 = 16'h2279; // 0x38be
	13'h1c60: q1 = 16'h0001; // 0x38c0
	13'h1c61: q1 = 16'h7eb2; // 0x38c2
	13'h1c62: q1 = 16'hd069; // 0x38c4
	13'h1c63: q1 = 16'h0004; // 0x38c6
	13'h1c64: q1 = 16'h3d40; // 0x38c8
	13'h1c65: q1 = 16'hfffc; // 0x38ca
	13'h1c66: q1 = 16'h302e; // 0x38cc
	13'h1c67: q1 = 16'hfffe; // 0x38ce
	13'h1c68: q1 = 16'h9079; // 0x38d0
	13'h1c69: q1 = 16'h0001; // 0x38d2
	13'h1c6a: q1 = 16'h861c; // 0x38d4
	13'h1c6b: q1 = 16'h33c0; // 0x38d6
	13'h1c6c: q1 = 16'h0001; // 0x38d8
	13'h1c6d: q1 = 16'h8622; // 0x38da
	13'h1c6e: q1 = 16'h3039; // 0x38dc
	13'h1c6f: q1 = 16'h0001; // 0x38de
	13'h1c70: q1 = 16'h8626; // 0x38e0
	13'h1c71: q1 = 16'h906e; // 0x38e2
	13'h1c72: q1 = 16'hfffc; // 0x38e4
	13'h1c73: q1 = 16'h33c0; // 0x38e6
	13'h1c74: q1 = 16'h0001; // 0x38e8
	13'h1c75: q1 = 16'h8624; // 0x38ea
	13'h1c76: q1 = 16'h4a9f; // 0x38ec
	13'h1c77: q1 = 16'h4cdf; // 0x38ee
	13'h1c78: q1 = 16'h2080; // 0x38f0
	13'h1c79: q1 = 16'h4e5e; // 0x38f2
	13'h1c7a: q1 = 16'h4e75; // 0x38f4
	13'h1c7b: q1 = 16'h4e56; // 0x38f6
	13'h1c7c: q1 = 16'h0000; // 0x38f8
	13'h1c7d: q1 = 16'h48e7; // 0x38fa
	13'h1c7e: q1 = 16'h1f1c; // 0x38fc
	13'h1c7f: q1 = 16'h2a6e; // 0x38fe
	13'h1c80: q1 = 16'h0008; // 0x3900
	13'h1c81: q1 = 16'h3e2e; // 0x3902
	13'h1c82: q1 = 16'h000c; // 0x3904
	13'h1c83: q1 = 16'hbe7c; // 0x3906
	13'h1c84: q1 = 16'h003c; // 0x3908
	13'h1c85: q1 = 16'h6e1c; // 0x390a
	13'h1c86: q1 = 16'h287c; // 0x390c
	13'h1c87: q1 = 16'h0000; // 0x390e
	13'h1c88: q1 = 16'he0e0; // 0x3910
	13'h1c89: q1 = 16'h3007; // 0x3912
	13'h1c8a: q1 = 16'he740; // 0x3914
	13'h1c8b: q1 = 16'h48c0; // 0x3916
	13'h1c8c: q1 = 16'hd9c0; // 0x3918
	13'h1c8d: q1 = 16'h3039; // 0x391a
	13'h1c8e: q1 = 16'h0001; // 0x391c
	13'h1c8f: q1 = 16'h758c; // 0x391e
	13'h1c90: q1 = 16'he340; // 0x3920
	13'h1c91: q1 = 16'h48c0; // 0x3922
	13'h1c92: q1 = 16'hd9c0; // 0x3924
	13'h1c93: q1 = 16'h6012; // 0x3926
	13'h1c94: q1 = 16'h287c; // 0x3928
	13'h1c95: q1 = 16'h0000; // 0x392a
	13'h1c96: q1 = 16'he2c8; // 0x392c
	13'h1c97: q1 = 16'h3007; // 0x392e
	13'h1c98: q1 = 16'hd07c; // 0x3930
	13'h1c99: q1 = 16'hffc3; // 0x3932
	13'h1c9a: q1 = 16'he340; // 0x3934
	13'h1c9b: q1 = 16'h48c0; // 0x3936
	13'h1c9c: q1 = 16'hd9c0; // 0x3938
	13'h1c9d: q1 = 16'h267c; // 0x393a
	13'h1c9e: q1 = 16'h0000; // 0x393c
	13'h1c9f: q1 = 16'he3b8; // 0x393e
	13'h1ca0: q1 = 16'h3014; // 0x3940
	13'h1ca1: q1 = 16'h48c0; // 0x3942
	13'h1ca2: q1 = 16'hd7c0; // 0x3944
	13'h1ca3: q1 = 16'h7803; // 0x3946
	13'h1ca4: q1 = 16'hb87c; // 0x3948
	13'h1ca5: q1 = 16'h0003; // 0x394a
	13'h1ca6: q1 = 16'h662e; // 0x394c
	13'h1ca7: q1 = 16'h101b; // 0x394e
	13'h1ca8: q1 = 16'h4880; // 0x3950
	13'h1ca9: q1 = 16'h48c0; // 0x3952
	13'h1caa: q1 = 16'h2c00; // 0x3954
	13'h1cab: q1 = 16'h4280; // 0x3956
	13'h1cac: q1 = 16'h7010; // 0x3958
	13'h1cad: q1 = 16'he1a6; // 0x395a
	13'h1cae: q1 = 16'h101b; // 0x395c
	13'h1caf: q1 = 16'h4880; // 0x395e
	13'h1cb0: q1 = 16'he140; // 0x3960
	13'h1cb1: q1 = 16'h48c0; // 0x3962
	13'h1cb2: q1 = 16'hc0b9; // 0x3964
	13'h1cb3: q1 = 16'h0000; // 0x3966
	13'h1cb4: q1 = 16'he3b4; // 0x3968
	13'h1cb5: q1 = 16'h8c80; // 0x396a
	13'h1cb6: q1 = 16'h101b; // 0x396c
	13'h1cb7: q1 = 16'h4880; // 0x396e
	13'h1cb8: q1 = 16'hc07c; // 0x3970
	13'h1cb9: q1 = 16'h00ff; // 0x3972
	13'h1cba: q1 = 16'h48c0; // 0x3974
	13'h1cbb: q1 = 16'h8c80; // 0x3976
	13'h1cbc: q1 = 16'h4244; // 0x3978
	13'h1cbd: q1 = 16'h6004; // 0x397a
	13'h1cbe: q1 = 16'hed86; // 0x397c
	13'h1cbf: q1 = 16'h5244; // 0x397e
	13'h1cc0: q1 = 16'h2006; // 0x3980
	13'h1cc1: q1 = 16'h4281; // 0x3982
	13'h1cc2: q1 = 16'h7212; // 0x3984
	13'h1cc3: q1 = 16'he2a0; // 0x3986
	13'h1cc4: q1 = 16'hc0bc; // 0x3988
	13'h1cc5: q1 = 16'h0000; // 0x398a
	13'h1cc6: q1 = 16'h003f; // 0x398c
	13'h1cc7: q1 = 16'h3a00; // 0x398e
	13'h1cc8: q1 = 16'hba7c; // 0x3990
	13'h1cc9: q1 = 16'h003e; // 0x3992
	13'h1cca: q1 = 16'h670a; // 0x3994
	13'h1ccb: q1 = 16'h3005; // 0x3996
	13'h1ccc: q1 = 16'hd07c; // 0x3998
	13'h1ccd: q1 = 16'h0020; // 0x399a
	13'h1cce: q1 = 16'h1ac0; // 0x399c
	13'h1ccf: q1 = 16'h60a8; // 0x399e
	13'h1cd0: q1 = 16'h4215; // 0x39a0
	13'h1cd1: q1 = 16'h4a9f; // 0x39a2
	13'h1cd2: q1 = 16'h4cdf; // 0x39a4
	13'h1cd3: q1 = 16'h38f0; // 0x39a6
	13'h1cd4: q1 = 16'h4e5e; // 0x39a8
	13'h1cd5: q1 = 16'h4e75; // 0x39aa
	13'h1cd6: q1 = 16'h4e56; // 0x39ac
	13'h1cd7: q1 = 16'h0000; // 0x39ae
	13'h1cd8: q1 = 16'h48e7; // 0x39b0
	13'h1cd9: q1 = 16'h3f00; // 0x39b2
	13'h1cda: q1 = 16'h4243; // 0x39b4
	13'h1cdb: q1 = 16'h2e2e; // 0x39b6
	13'h1cdc: q1 = 16'h0008; // 0x39b8
	13'h1cdd: q1 = 16'h2c2e; // 0x39ba
	13'h1cde: q1 = 16'h000c; // 0x39bc
	13'h1cdf: q1 = 16'h4a86; // 0x39be
	13'h1ce0: q1 = 16'h6614; // 0x39c0
	13'h1ce1: q1 = 16'h23f9; // 0x39c2
	13'h1ce2: q1 = 16'h0000; // 0x39c4
	13'h1ce3: q1 = 16'hf316; // 0x39c6
	13'h1ce4: q1 = 16'h0001; // 0x39c8
	13'h1ce5: q1 = 16'h81f6; // 0x39ca
	13'h1ce6: q1 = 16'h2039; // 0x39cc
	13'h1ce7: q1 = 16'h0000; // 0x39ce
	13'h1ce8: q1 = 16'hf316; // 0x39d0
	13'h1ce9: q1 = 16'h6000; // 0x39d2
	13'h1cea: q1 = 16'h0072; // 0x39d4
	13'h1ceb: q1 = 16'h4a87; // 0x39d6
	13'h1cec: q1 = 16'h6c08; // 0x39d8
	13'h1ced: q1 = 16'h2007; // 0x39da
	13'h1cee: q1 = 16'h4480; // 0x39dc
	13'h1cef: q1 = 16'h2e00; // 0x39de
	13'h1cf0: q1 = 16'h5243; // 0x39e0
	13'h1cf1: q1 = 16'h4a86; // 0x39e2
	13'h1cf2: q1 = 16'h6c08; // 0x39e4
	13'h1cf3: q1 = 16'h2006; // 0x39e6
	13'h1cf4: q1 = 16'h4480; // 0x39e8
	13'h1cf5: q1 = 16'h2c00; // 0x39ea
	13'h1cf6: q1 = 16'h5243; // 0x39ec
	13'h1cf7: q1 = 16'hbc87; // 0x39ee
	13'h1cf8: q1 = 16'h6f0c; // 0x39f0
	13'h1cf9: q1 = 16'h23ee; // 0x39f2
	13'h1cfa: q1 = 16'h0008; // 0x39f4
	13'h1cfb: q1 = 16'h0001; // 0x39f6
	13'h1cfc: q1 = 16'h81f6; // 0x39f8
	13'h1cfd: q1 = 16'h7000; // 0x39fa
	13'h1cfe: q1 = 16'h6048; // 0x39fc
	13'h1cff: q1 = 16'hbe86; // 0x39fe
	13'h1d00: q1 = 16'h6606; // 0x3a00
	13'h1d01: q1 = 16'h7a01; // 0x3a02
	13'h1d02: q1 = 16'h4287; // 0x3a04
	13'h1d03: q1 = 16'h6020; // 0x3a06
	13'h1d04: q1 = 16'h7801; // 0x3a08
	13'h1d05: q1 = 16'hbe86; // 0x3a0a
	13'h1d06: q1 = 16'h6d06; // 0x3a0c
	13'h1d07: q1 = 16'he386; // 0x3a0e
	13'h1d08: q1 = 16'he384; // 0x3a10
	13'h1d09: q1 = 16'h60f6; // 0x3a12
	13'h1d0a: q1 = 16'h4285; // 0x3a14
	13'h1d0b: q1 = 16'h4a84; // 0x3a16
	13'h1d0c: q1 = 16'h670e; // 0x3a18
	13'h1d0d: q1 = 16'hbe86; // 0x3a1a
	13'h1d0e: q1 = 16'h6d04; // 0x3a1c
	13'h1d0f: q1 = 16'h8a84; // 0x3a1e
	13'h1d10: q1 = 16'h9e86; // 0x3a20
	13'h1d11: q1 = 16'he284; // 0x3a22
	13'h1d12: q1 = 16'he286; // 0x3a24
	13'h1d13: q1 = 16'h60ee; // 0x3a26
	13'h1d14: q1 = 16'hb67c; // 0x3a28
	13'h1d15: q1 = 16'h0001; // 0x3a2a
	13'h1d16: q1 = 16'h6610; // 0x3a2c
	13'h1d17: q1 = 16'h2007; // 0x3a2e
	13'h1d18: q1 = 16'h4480; // 0x3a30
	13'h1d19: q1 = 16'h23c0; // 0x3a32
	13'h1d1a: q1 = 16'h0001; // 0x3a34
	13'h1d1b: q1 = 16'h81f6; // 0x3a36
	13'h1d1c: q1 = 16'h2005; // 0x3a38
	13'h1d1d: q1 = 16'h4480; // 0x3a3a
	13'h1d1e: q1 = 16'h6008; // 0x3a3c
	13'h1d1f: q1 = 16'h23c7; // 0x3a3e
	13'h1d20: q1 = 16'h0001; // 0x3a40
	13'h1d21: q1 = 16'h81f6; // 0x3a42
	13'h1d22: q1 = 16'h2005; // 0x3a44
	13'h1d23: q1 = 16'h4a9f; // 0x3a46
	13'h1d24: q1 = 16'h4cdf; // 0x3a48
	13'h1d25: q1 = 16'h00f8; // 0x3a4a
	13'h1d26: q1 = 16'h4e5e; // 0x3a4c
	13'h1d27: q1 = 16'h4e75; // 0x3a4e
	13'h1d28: q1 = 16'h4e56; // 0x3a50
	13'h1d29: q1 = 16'hfffc; // 0x3a52
	13'h1d2a: q1 = 16'h4242; // 0x3a54
	13'h1d2b: q1 = 16'h4aae; // 0x3a56
	13'h1d2c: q1 = 16'h0008; // 0x3a58
	13'h1d2d: q1 = 16'h6c06; // 0x3a5a
	13'h1d2e: q1 = 16'h44ae; // 0x3a5c
	13'h1d2f: q1 = 16'h0008; // 0x3a5e
	13'h1d30: q1 = 16'h5242; // 0x3a60
	13'h1d31: q1 = 16'h4aae; // 0x3a62
	13'h1d32: q1 = 16'h000c; // 0x3a64
	13'h1d33: q1 = 16'h6c06; // 0x3a66
	13'h1d34: q1 = 16'h44ae; // 0x3a68
	13'h1d35: q1 = 16'h000c; // 0x3a6a
	13'h1d36: q1 = 16'h5242; // 0x3a6c
	13'h1d37: q1 = 16'h302e; // 0x3a6e
	13'h1d38: q1 = 16'h000a; // 0x3a70
	13'h1d39: q1 = 16'hc0ee; // 0x3a72
	13'h1d3a: q1 = 16'h000e; // 0x3a74
	13'h1d3b: q1 = 16'h2d40; // 0x3a76
	13'h1d3c: q1 = 16'hfffc; // 0x3a78
	13'h1d3d: q1 = 16'h302e; // 0x3a7a
	13'h1d3e: q1 = 16'h0008; // 0x3a7c
	13'h1d3f: q1 = 16'hc0ee; // 0x3a7e
	13'h1d40: q1 = 16'h000e; // 0x3a80
	13'h1d41: q1 = 16'h322e; // 0x3a82
	13'h1d42: q1 = 16'h000c; // 0x3a84
	13'h1d43: q1 = 16'hc2ee; // 0x3a86
	13'h1d44: q1 = 16'h000a; // 0x3a88
	13'h1d45: q1 = 16'hd041; // 0x3a8a
	13'h1d46: q1 = 16'hd06e; // 0x3a8c
	13'h1d47: q1 = 16'hfffc; // 0x3a8e
	13'h1d48: q1 = 16'h3d40; // 0x3a90
	13'h1d49: q1 = 16'hfffc; // 0x3a92
	13'h1d4a: q1 = 16'h202e; // 0x3a94
	13'h1d4b: q1 = 16'hfffc; // 0x3a96
	13'h1d4c: q1 = 16'h0802; // 0x3a98
	13'h1d4d: q1 = 16'h0000; // 0x3a9a
	13'h1d4e: q1 = 16'h6702; // 0x3a9c
	13'h1d4f: q1 = 16'h4480; // 0x3a9e
	13'h1d50: q1 = 16'h4e5e; // 0x3aa0
	13'h1d51: q1 = 16'h4e75; // 0x3aa2
	13'h1d52: q1 = 16'h4e56; // 0x3aa4
	13'h1d53: q1 = 16'hfff6; // 0x3aa6
	13'h1d54: q1 = 16'h48e7; // 0x3aa8
	13'h1d55: q1 = 16'h3f04; // 0x3aaa
	13'h1d56: q1 = 16'h33fc; // 0x3aac
	13'h1d57: q1 = 16'h0001; // 0x3aae
	13'h1d58: q1 = 16'h0001; // 0x3ab0
	13'h1d59: q1 = 16'h7f1c; // 0x3ab2
	13'h1d5a: q1 = 16'h4279; // 0x3ab4
	13'h1d5b: q1 = 16'h0001; // 0x3ab6
	13'h1d5c: q1 = 16'h7f1e; // 0x3ab8
	13'h1d5d: q1 = 16'h4247; // 0x3aba
	13'h1d5e: q1 = 16'hbe7c; // 0x3abc
	13'h1d5f: q1 = 16'h0020; // 0x3abe
	13'h1d60: q1 = 16'h6c00; // 0x3ac0
	13'h1d61: q1 = 16'h0118; // 0x3ac2
	13'h1d62: q1 = 16'h7c1f; // 0x3ac4
	13'h1d63: q1 = 16'hbc7c; // 0x3ac6
	13'h1d64: q1 = 16'h0019; // 0x3ac8
	13'h1d65: q1 = 16'h6d00; // 0x3aca
	13'h1d66: q1 = 16'h0108; // 0x3acc
	13'h1d67: q1 = 16'h3007; // 0x3ace
	13'h1d68: q1 = 16'h48c0; // 0x3ad0
	13'h1d69: q1 = 16'hd0bc; // 0x3ad2
	13'h1d6a: q1 = 16'h0000; // 0x3ad4
	13'h1d6b: q1 = 16'hf356; // 0x3ad6
	13'h1d6c: q1 = 16'h2040; // 0x3ad8
	13'h1d6d: q1 = 16'h1010; // 0x3ada
	13'h1d6e: q1 = 16'h4880; // 0x3adc
	13'h1d6f: q1 = 16'h4281; // 0x3ade
	13'h1d70: q1 = 16'h3206; // 0x3ae0
	13'h1d71: q1 = 16'hd27c; // 0x3ae2
	13'h1d72: q1 = 16'hffe7; // 0x3ae4
	13'h1d73: q1 = 16'he260; // 0x3ae6
	13'h1d74: q1 = 16'hc07c; // 0x3ae8
	13'h1d75: q1 = 16'h0001; // 0x3aea
	13'h1d76: q1 = 16'h6700; // 0x3aec
	13'h1d77: q1 = 16'h00e0; // 0x3aee
	13'h1d78: q1 = 16'h4243; // 0x3af0
	13'h1d79: q1 = 16'h23fc; // 0x3af2
	13'h1d7a: q1 = 16'h0000; // 0x3af4
	13'h1d7b: q1 = 16'h0002; // 0x3af6
	13'h1d7c: q1 = 16'h0001; // 0x3af8
	13'h1d7d: q1 = 16'h7fc2; // 0x3afa
	13'h1d7e: q1 = 16'h3ebc; // 0x3afc
	13'h1d7f: q1 = 16'h7880; // 0x3afe
	13'h1d80: q1 = 16'h3f3c; // 0x3b00
	13'h1d81: q1 = 16'h0080; // 0x3b02
	13'h1d82: q1 = 16'h4eb9; // 0x3b04
	13'h1d83: q1 = 16'h0000; // 0x3b06
	13'h1d84: q1 = 16'h8e6c; // 0x3b08
	13'h1d85: q1 = 16'h4a5f; // 0x3b0a
	13'h1d86: q1 = 16'h3a00; // 0x3b0c
	13'h1d87: q1 = 16'h383c; // 0x3b0e
	13'h1d88: q1 = 16'h1280; // 0x3b10
	13'h1d89: q1 = 16'h3ebc; // 0x3b12
	13'h1d8a: q1 = 16'h0005; // 0x3b14
	13'h1d8b: q1 = 16'h3f3c; // 0x3b16
	13'h1d8c: q1 = 16'h0001; // 0x3b18
	13'h1d8d: q1 = 16'h4eb9; // 0x3b1a
	13'h1d8e: q1 = 16'h0000; // 0x3b1c
	13'h1d8f: q1 = 16'h8e6c; // 0x3b1e
	13'h1d90: q1 = 16'h4a5f; // 0x3b20
	13'h1d91: q1 = 16'h3d40; // 0x3b22
	13'h1d92: q1 = 16'hfff6; // 0x3b24
	13'h1d93: q1 = 16'h3007; // 0x3b26
	13'h1d94: q1 = 16'h4281; // 0x3b28
	13'h1d95: q1 = 16'h720a; // 0x3b2a
	13'h1d96: q1 = 16'he360; // 0x3b2c
	13'h1d97: q1 = 16'hd07c; // 0x3b2e
	13'h1d98: q1 = 16'hfe00; // 0x3b30
	13'h1d99: q1 = 16'h3d40; // 0x3b32
	13'h1d9a: q1 = 16'hfffa; // 0x3b34
	13'h1d9b: q1 = 16'h3006; // 0x3b36
	13'h1d9c: q1 = 16'h4281; // 0x3b38
	13'h1d9d: q1 = 16'h720a; // 0x3b3a
	13'h1d9e: q1 = 16'he360; // 0x3b3c
	13'h1d9f: q1 = 16'hd07c; // 0x3b3e
	13'h1da0: q1 = 16'hfe00; // 0x3b40
	13'h1da1: q1 = 16'h3d40; // 0x3b42
	13'h1da2: q1 = 16'hfff8; // 0x3b44
	13'h1da3: q1 = 16'h3e84; // 0x3b46
	13'h1da4: q1 = 16'h3f05; // 0x3b48
	13'h1da5: q1 = 16'h3f2e; // 0x3b4a
	13'h1da6: q1 = 16'hfff6; // 0x3b4c
	13'h1da7: q1 = 16'h4eb9; // 0x3b4e
	13'h1da8: q1 = 16'h0000; // 0x3b50
	13'h1da9: q1 = 16'h38d8; // 0x3b52
	13'h1daa: q1 = 16'h4a9f; // 0x3b54
	13'h1dab: q1 = 16'h2a40; // 0x3b56
	13'h1dac: q1 = 16'h200d; // 0x3b58
	13'h1dad: q1 = 16'h6752; // 0x3b5a
	13'h1dae: q1 = 16'h302e; // 0x3b5c
	13'h1daf: q1 = 16'hfffa; // 0x3b5e
	13'h1db0: q1 = 16'h9045; // 0x3b60
	13'h1db1: q1 = 16'h3d40; // 0x3b62
	13'h1db2: q1 = 16'hfffe; // 0x3b64
	13'h1db3: q1 = 16'h302e; // 0x3b66
	13'h1db4: q1 = 16'hfff8; // 0x3b68
	13'h1db5: q1 = 16'h9044; // 0x3b6a
	13'h1db6: q1 = 16'h3d40; // 0x3b6c
	13'h1db7: q1 = 16'hfffc; // 0x3b6e
	13'h1db8: q1 = 16'h200e; // 0x3b70
	13'h1db9: q1 = 16'hd0bc; // 0x3b72
	13'h1dba: q1 = 16'hffff; // 0x3b74
	13'h1dbb: q1 = 16'hfffc; // 0x3b76
	13'h1dbc: q1 = 16'h2e80; // 0x3b78
	13'h1dbd: q1 = 16'h200e; // 0x3b7a
	13'h1dbe: q1 = 16'hd0bc; // 0x3b7c
	13'h1dbf: q1 = 16'hffff; // 0x3b7e
	13'h1dc0: q1 = 16'hfffe; // 0x3b80
	13'h1dc1: q1 = 16'h2f00; // 0x3b82
	13'h1dc2: q1 = 16'h3f3c; // 0x3b84
	13'h1dc3: q1 = 16'h0600; // 0x3b86
	13'h1dc4: q1 = 16'h4eb9; // 0x3b88
	13'h1dc5: q1 = 16'h0000; // 0x3b8a
	13'h1dc6: q1 = 16'h09bc; // 0x3b8c
	13'h1dc7: q1 = 16'h5c4f; // 0x3b8e
	13'h1dc8: q1 = 16'h3eae; // 0x3b90
	13'h1dc9: q1 = 16'hfff8; // 0x3b92
	13'h1dca: q1 = 16'h3f2e; // 0x3b94
	13'h1dcb: q1 = 16'hfffa; // 0x3b96
	13'h1dcc: q1 = 16'h3f2e; // 0x3b98
	13'h1dcd: q1 = 16'hfffc; // 0x3b9a
	13'h1dce: q1 = 16'h3f2e; // 0x3b9c
	13'h1dcf: q1 = 16'hfffe; // 0x3b9e
	13'h1dd0: q1 = 16'h2f0d; // 0x3ba0
	13'h1dd1: q1 = 16'h4eb9; // 0x3ba2
	13'h1dd2: q1 = 16'h0000; // 0x3ba4
	13'h1dd3: q1 = 16'h3988; // 0x3ba6
	13'h1dd4: q1 = 16'hdefc; // 0x3ba8
	13'h1dd5: q1 = 16'h000a; // 0x3baa
	13'h1dd6: q1 = 16'h5243; // 0x3bac
	13'h1dd7: q1 = 16'h4eb9; // 0x3bae
	13'h1dd8: q1 = 16'h0000; // 0x3bb0
	13'h1dd9: q1 = 16'h2fb4; // 0x3bb2
	13'h1dda: q1 = 16'h4ab9; // 0x3bb4
	13'h1ddb: q1 = 16'h0001; // 0x3bb6
	13'h1ddc: q1 = 16'h7fc2; // 0x3bb8
	13'h1ddd: q1 = 16'h670a; // 0x3bba
	13'h1dde: q1 = 16'h4a79; // 0x3bbc
	13'h1ddf: q1 = 16'h0001; // 0x3bbe
	13'h1de0: q1 = 16'h7594; // 0x3bc0
	13'h1de1: q1 = 16'h6616; // 0x3bc2
	13'h1de2: q1 = 16'h60ee; // 0x3bc4
	13'h1de3: q1 = 16'h4a43; // 0x3bc6
	13'h1de4: q1 = 16'h6e04; // 0x3bc8
	13'h1de5: q1 = 16'h6000; // 0x3bca
	13'h1de6: q1 = 16'hff26; // 0x3bcc
	13'h1de7: q1 = 16'h5346; // 0x3bce
	13'h1de8: q1 = 16'h6000; // 0x3bd0
	13'h1de9: q1 = 16'hfef4; // 0x3bd2
	13'h1dea: q1 = 16'h5247; // 0x3bd4
	13'h1deb: q1 = 16'h6000; // 0x3bd6
	13'h1dec: q1 = 16'hfee4; // 0x3bd8
	13'h1ded: q1 = 16'h4279; // 0x3bda
	13'h1dee: q1 = 16'h0001; // 0x3bdc
	13'h1def: q1 = 16'h7f1c; // 0x3bde
	13'h1df0: q1 = 16'h4a9f; // 0x3be0
	13'h1df1: q1 = 16'h4cdf; // 0x3be2
	13'h1df2: q1 = 16'h20f8; // 0x3be4
	13'h1df3: q1 = 16'h4e5e; // 0x3be6
	13'h1df4: q1 = 16'h4e75; // 0x3be8
	13'h1df5: q1 = 16'h4e56; // 0x3bea
	13'h1df6: q1 = 16'hfffc; // 0x3bec
	13'h1df7: q1 = 16'h4eb9; // 0x3bee
	13'h1df8: q1 = 16'h0000; // 0x3bf0
	13'h1df9: q1 = 16'h6316; // 0x3bf2
	13'h1dfa: q1 = 16'h4279; // 0x3bf4
	13'h1dfb: q1 = 16'h0001; // 0x3bf6
	13'h1dfc: q1 = 16'h867a; // 0x3bf8
	13'h1dfd: q1 = 16'h33fc; // 0x3bfa
	13'h1dfe: q1 = 16'h0001; // 0x3bfc
	13'h1dff: q1 = 16'h0001; // 0x3bfe
	13'h1e00: q1 = 16'h7fc6; // 0x3c00
	13'h1e01: q1 = 16'h4eb9; // 0x3c02
	13'h1e02: q1 = 16'h0000; // 0x3c04
	13'h1e03: q1 = 16'h2304; // 0x3c06
	13'h1e04: q1 = 16'h3ebc; // 0x3c08
	13'h1e05: q1 = 16'h0004; // 0x3c0a
	13'h1e06: q1 = 16'h4eb9; // 0x3c0c
	13'h1e07: q1 = 16'h0000; // 0x3c0e
	13'h1e08: q1 = 16'h0aaa; // 0x3c10
	13'h1e09: q1 = 16'h4a79; // 0x3c12
	13'h1e0a: q1 = 16'h0001; // 0x3c14
	13'h1e0b: q1 = 16'h7f5e; // 0x3c16
	13'h1e0c: q1 = 16'h6652; // 0x3c18
	13'h1e0d: q1 = 16'h3ebc; // 0x3c1a
	13'h1e0e: q1 = 16'h000f; // 0x3c1c
	13'h1e0f: q1 = 16'h4eb9; // 0x3c1e
	13'h1e10: q1 = 16'h0000; // 0x3c20
	13'h1e11: q1 = 16'h0aaa; // 0x3c22
	13'h1e12: q1 = 16'h4a79; // 0x3c24
	13'h1e13: q1 = 16'h0001; // 0x3c26
	13'h1e14: q1 = 16'h7f5e; // 0x3c28
	13'h1e15: q1 = 16'h6640; // 0x3c2a
	13'h1e16: q1 = 16'h4a79; // 0x3c2c
	13'h1e17: q1 = 16'h0001; // 0x3c2e
	13'h1e18: q1 = 16'h7594; // 0x3c30
	13'h1e19: q1 = 16'h6606; // 0x3c32
	13'h1e1a: q1 = 16'h4eb9; // 0x3c34
	13'h1e1b: q1 = 16'h0000; // 0x3c36
	13'h1e1c: q1 = 16'h6d02; // 0x3c38
	13'h1e1d: q1 = 16'h4a79; // 0x3c3a
	13'h1e1e: q1 = 16'h0001; // 0x3c3c
	13'h1e1f: q1 = 16'h7f5e; // 0x3c3e
	13'h1e20: q1 = 16'h662a; // 0x3c40
	13'h1e21: q1 = 16'h3ebc; // 0x3c42
	13'h1e22: q1 = 16'h0020; // 0x3c44
	13'h1e23: q1 = 16'h4eb9; // 0x3c46
	13'h1e24: q1 = 16'h0000; // 0x3c48
	13'h1e25: q1 = 16'h0aaa; // 0x3c4a
	13'h1e26: q1 = 16'h4a79; // 0x3c4c
	13'h1e27: q1 = 16'h0001; // 0x3c4e
	13'h1e28: q1 = 16'h7f5e; // 0x3c50
	13'h1e29: q1 = 16'h6618; // 0x3c52
	13'h1e2a: q1 = 16'h4a79; // 0x3c54
	13'h1e2b: q1 = 16'h0001; // 0x3c56
	13'h1e2c: q1 = 16'h7594; // 0x3c58
	13'h1e2d: q1 = 16'h6606; // 0x3c5a
	13'h1e2e: q1 = 16'h4eb9; // 0x3c5c
	13'h1e2f: q1 = 16'h0000; // 0x3c5e
	13'h1e30: q1 = 16'hb49a; // 0x3c60
	13'h1e31: q1 = 16'h4a79; // 0x3c62
	13'h1e32: q1 = 16'h0001; // 0x3c64
	13'h1e33: q1 = 16'h7f5e; // 0x3c66
	13'h1e34: q1 = 16'h6602; // 0x3c68
	13'h1e35: q1 = 16'h6096; // 0x3c6a
	13'h1e36: q1 = 16'h4ab9; // 0x3c6c
	13'h1e37: q1 = 16'h0001; // 0x3c6e
	13'h1e38: q1 = 16'h7fac; // 0x3c70
	13'h1e39: q1 = 16'h6614; // 0x3c72
	13'h1e3a: q1 = 16'h33fc; // 0x3c74
	13'h1e3b: q1 = 16'h0001; // 0x3c76
	13'h1e3c: q1 = 16'h0001; // 0x3c78
	13'h1e3d: q1 = 16'h7eb6; // 0x3c7a
	13'h1e3e: q1 = 16'h4279; // 0x3c7c
	13'h1e3f: q1 = 16'h0001; // 0x3c7e
	13'h1e40: q1 = 16'h8644; // 0x3c80
	13'h1e41: q1 = 16'h4279; // 0x3c82
	13'h1e42: q1 = 16'h0001; // 0x3c84
	13'h1e43: q1 = 16'h866a; // 0x3c86
	13'h1e44: q1 = 16'h33fc; // 0x3c88
	13'h1e45: q1 = 16'h0001; // 0x3c8a
	13'h1e46: q1 = 16'h0001; // 0x3c8c
	13'h1e47: q1 = 16'h867a; // 0x3c8e
	13'h1e48: q1 = 16'h4279; // 0x3c90
	13'h1e49: q1 = 16'h0001; // 0x3c92
	13'h1e4a: q1 = 16'h7fc6; // 0x3c94
	13'h1e4b: q1 = 16'h4eb9; // 0x3c96
	13'h1e4c: q1 = 16'h0000; // 0x3c98
	13'h1e4d: q1 = 16'h44ac; // 0x3c9a
	13'h1e4e: q1 = 16'h4eb9; // 0x3c9c
	13'h1e4f: q1 = 16'h0000; // 0x3c9e
	13'h1e50: q1 = 16'h827e; // 0x3ca0
	13'h1e51: q1 = 16'h0c79; // 0x3ca2
	13'h1e52: q1 = 16'h0001; // 0x3ca4
	13'h1e53: q1 = 16'h0001; // 0x3ca6
	13'h1e54: q1 = 16'h87dc; // 0x3ca8
	13'h1e55: q1 = 16'h660c; // 0x3caa
	13'h1e56: q1 = 16'h33f9; // 0x3cac
	13'h1e57: q1 = 16'h0001; // 0x3cae
	13'h1e58: q1 = 16'h8628; // 0x3cb0
	13'h1e59: q1 = 16'h0001; // 0x3cb2
	13'h1e5a: q1 = 16'h7eb6; // 0x3cb4
	13'h1e5b: q1 = 16'h6024; // 0x3cb6
	13'h1e5c: q1 = 16'h3039; // 0x3cb8
	13'h1e5d: q1 = 16'h0001; // 0x3cba
	13'h1e5e: q1 = 16'h8628; // 0x3cbc
	13'h1e5f: q1 = 16'hb079; // 0x3cbe
	13'h1e60: q1 = 16'h0001; // 0x3cc0
	13'h1e61: q1 = 16'h864e; // 0x3cc2
	13'h1e62: q1 = 16'h6f0c; // 0x3cc4
	13'h1e63: q1 = 16'h33f9; // 0x3cc6
	13'h1e64: q1 = 16'h0001; // 0x3cc8
	13'h1e65: q1 = 16'h8628; // 0x3cca
	13'h1e66: q1 = 16'h0001; // 0x3ccc
	13'h1e67: q1 = 16'h7eb6; // 0x3cce
	13'h1e68: q1 = 16'h600a; // 0x3cd0
	13'h1e69: q1 = 16'h33f9; // 0x3cd2
	13'h1e6a: q1 = 16'h0001; // 0x3cd4
	13'h1e6b: q1 = 16'h864e; // 0x3cd6
	13'h1e6c: q1 = 16'h0001; // 0x3cd8
	13'h1e6d: q1 = 16'h7eb6; // 0x3cda
	13'h1e6e: q1 = 16'h0c79; // 0x3cdc
	13'h1e6f: q1 = 16'h0001; // 0x3cde
	13'h1e70: q1 = 16'h0001; // 0x3ce0
	13'h1e71: q1 = 16'h7eb6; // 0x3ce2
	13'h1e72: q1 = 16'h660e; // 0x3ce4
	13'h1e73: q1 = 16'h4279; // 0x3ce6
	13'h1e74: q1 = 16'h0001; // 0x3ce8
	13'h1e75: q1 = 16'h8644; // 0x3cea
	13'h1e76: q1 = 16'h4279; // 0x3cec
	13'h1e77: q1 = 16'h0001; // 0x3cee
	13'h1e78: q1 = 16'h866a; // 0x3cf0
	13'h1e79: q1 = 16'h6010; // 0x3cf2
	13'h1e7a: q1 = 16'h33fc; // 0x3cf4
	13'h1e7b: q1 = 16'h0001; // 0x3cf6
	13'h1e7c: q1 = 16'h0001; // 0x3cf8
	13'h1e7d: q1 = 16'h8644; // 0x3cfa
	13'h1e7e: q1 = 16'h33fc; // 0x3cfc
	13'h1e7f: q1 = 16'h0001; // 0x3cfe
	13'h1e80: q1 = 16'h0001; // 0x3d00
	13'h1e81: q1 = 16'h866a; // 0x3d02
	13'h1e82: q1 = 16'h4279; // 0x3d04
	13'h1e83: q1 = 16'h0001; // 0x3d06
	13'h1e84: q1 = 16'h867a; // 0x3d08
	13'h1e85: q1 = 16'h3eb9; // 0x3d0a
	13'h1e86: q1 = 16'h0001; // 0x3d0c
	13'h1e87: q1 = 16'h8054; // 0x3d0e
	13'h1e88: q1 = 16'h4eb9; // 0x3d10
	13'h1e89: q1 = 16'h0000; // 0x3d12
	13'h1e8a: q1 = 16'h64bc; // 0x3d14
	13'h1e8b: q1 = 16'h4a79; // 0x3d16
	13'h1e8c: q1 = 16'h0001; // 0x3d18
	13'h1e8d: q1 = 16'h7f5e; // 0x3d1a
	13'h1e8e: q1 = 16'h6600; // 0x3d1c
	13'h1e8f: q1 = 16'hff6a; // 0x3d1e
	13'h1e90: q1 = 16'h0c79; // 0x3d20
	13'h1e91: q1 = 16'h0002; // 0x3d22
	13'h1e92: q1 = 16'h0001; // 0x3d24
	13'h1e93: q1 = 16'h87dc; // 0x3d26
	13'h1e94: q1 = 16'h6612; // 0x3d28
	13'h1e95: q1 = 16'h3ebc; // 0x3d2a
	13'h1e96: q1 = 16'h0001; // 0x3d2c
	13'h1e97: q1 = 16'h3039; // 0x3d2e
	13'h1e98: q1 = 16'h0001; // 0x3d30
	13'h1e99: q1 = 16'h8054; // 0x3d32
	13'h1e9a: q1 = 16'h9157; // 0x3d34
	13'h1e9b: q1 = 16'h4eb9; // 0x3d36
	13'h1e9c: q1 = 16'h0000; // 0x3d38
	13'h1e9d: q1 = 16'h64bc; // 0x3d3a
	13'h1e9e: q1 = 16'h4eb9; // 0x3d3c
	13'h1e9f: q1 = 16'h0000; // 0x3d3e
	13'h1ea0: q1 = 16'h0226; // 0x3d40
	13'h1ea1: q1 = 16'h4a79; // 0x3d42
	13'h1ea2: q1 = 16'h0001; // 0x3d44
	13'h1ea3: q1 = 16'h758e; // 0x3d46
	13'h1ea4: q1 = 16'h670c; // 0x3d48
	13'h1ea5: q1 = 16'h4279; // 0x3d4a
	13'h1ea6: q1 = 16'h0001; // 0x3d4c
	13'h1ea7: q1 = 16'h7fa6; // 0x3d4e
	13'h1ea8: q1 = 16'h4279; // 0x3d50
	13'h1ea9: q1 = 16'h0001; // 0x3d52
	13'h1eaa: q1 = 16'h8052; // 0x3d54
	13'h1eab: q1 = 16'h4a79; // 0x3d56
	13'h1eac: q1 = 16'h0001; // 0x3d58
	13'h1ead: q1 = 16'h7f5e; // 0x3d5a
	13'h1eae: q1 = 16'h6600; // 0x3d5c
	13'h1eaf: q1 = 16'hff2a; // 0x3d5e
	13'h1eb0: q1 = 16'h4eb9; // 0x3d60
	13'h1eb1: q1 = 16'h0000; // 0x3d62
	13'h1eb2: q1 = 16'hb49a; // 0x3d64
	13'h1eb3: q1 = 16'h4a79; // 0x3d66
	13'h1eb4: q1 = 16'h0001; // 0x3d68
	13'h1eb5: q1 = 16'h7f5e; // 0x3d6a
	13'h1eb6: q1 = 16'h6600; // 0x3d6c
	13'h1eb7: q1 = 16'hff1a; // 0x3d6e
	13'h1eb8: q1 = 16'h23fc; // 0x3d70
	13'h1eb9: q1 = 16'h0000; // 0x3d72
	13'h1eba: q1 = 16'h0384; // 0x3d74
	13'h1ebb: q1 = 16'h0001; // 0x3d76
	13'h1ebc: q1 = 16'h7fac; // 0x3d78
	13'h1ebd: q1 = 16'h6004; // 0x3d7a
	13'h1ebe: q1 = 16'h6000; // 0x3d7c
	13'h1ebf: q1 = 16'hff0a; // 0x3d7e
	13'h1ec0: q1 = 16'h6000; // 0x3d80
	13'h1ec1: q1 = 16'hfe72; // 0x3d82
	13'h1ec2: q1 = 16'h4e5e; // 0x3d84
	13'h1ec3: q1 = 16'h4e75; // 0x3d86
	13'h1ec4: q1 = 16'h4e56; // 0x3d88
	13'h1ec5: q1 = 16'h0000; // 0x3d8a
	13'h1ec6: q1 = 16'h2f03; // 0x3d8c
	13'h1ec7: q1 = 16'h302e; // 0x3d8e
	13'h1ec8: q1 = 16'h0008; // 0x3d90
	13'h1ec9: q1 = 16'h207c; // 0x3d92
	13'h1eca: q1 = 16'h0000; // 0x3d94
	13'h1ecb: q1 = 16'hf4b6; // 0x3d96
	13'h1ecc: q1 = 16'hb058; // 0x3d98
	13'h1ecd: q1 = 16'h6cfc; // 0x3d9a
	13'h1ece: q1 = 16'h4281; // 0x3d9c
	13'h1ecf: q1 = 16'h3228; // 0x3d9e
	13'h1ed0: q1 = 16'h000e; // 0x3da0
	13'h1ed1: q1 = 16'he189; // 0x3da2
	13'h1ed2: q1 = 16'he389; // 0x3da4
	13'h1ed3: q1 = 16'h82c0; // 0x3da6
	13'h1ed4: q1 = 16'h3601; // 0x3da8
	13'h1ed5: q1 = 16'h4843; // 0x3daa
	13'h1ed6: q1 = 16'h4241; // 0x3dac
	13'h1ed7: q1 = 16'h82c0; // 0x3dae
	13'h1ed8: q1 = 16'h3601; // 0x3db0
	13'h1ed9: q1 = 16'h2408; // 0x3db2
	13'h1eda: q1 = 16'h94bc; // 0x3db4
	13'h1edb: q1 = 16'h0000; // 0x3db6
	13'h1edc: q1 = 16'hf4b8; // 0x3db8
	13'h1edd: q1 = 16'he38a; // 0x3dba
	13'h1ede: q1 = 16'hd4bc; // 0x3dbc
	13'h1edf: q1 = 16'h0000; // 0x3dbe
	13'h1ee0: q1 = 16'hf4d6; // 0x3dc0
	13'h1ee1: q1 = 16'h2042; // 0x3dc2
	13'h1ee2: q1 = 16'h2f10; // 0x3dc4
	13'h1ee3: q1 = 16'h4eb9; // 0x3dc6
	13'h1ee4: q1 = 16'h0000; // 0x3dc8
	13'h1ee5: q1 = 16'h7ff8; // 0x3dca
	13'h1ee6: q1 = 16'h588f; // 0x3dcc
	13'h1ee7: q1 = 16'h2143; // 0x3dce
	13'h1ee8: q1 = 16'h0000; // 0x3dd0
	13'h1ee9: q1 = 16'h261f; // 0x3dd2
	13'h1eea: q1 = 16'h4e5e; // 0x3dd4
	13'h1eeb: q1 = 16'h4e75; // 0x3dd6
	13'h1eec: q1 = 16'h3039; // 0x3dd8
	13'h1eed: q1 = 16'h0001; // 0x3dda
	13'h1eee: q1 = 16'h758a; // 0x3ddc
	13'h1eef: q1 = 16'h4640; // 0x3dde
	13'h1ef0: q1 = 16'hc079; // 0x3de0
	13'h1ef1: q1 = 16'h0001; // 0x3de2
	13'h1ef2: q1 = 16'h7fc6; // 0x3de4
	13'h1ef3: q1 = 16'h6704; // 0x3de6
	13'h1ef4: q1 = 16'h4240; // 0x3de8
	13'h1ef5: q1 = 16'h4e75; // 0x3dea
	13'h1ef6: q1 = 16'h4e56; // 0x3dec
	13'h1ef7: q1 = 16'hfffc; // 0x3dee
	13'h1ef8: q1 = 16'h4eb9; // 0x3df0
	13'h1ef9: q1 = 16'h0000; // 0x3df2
	13'h1efa: q1 = 16'h01de; // 0x3df4
	13'h1efb: q1 = 16'h2eae; // 0x3df6
	13'h1efc: q1 = 16'h0008; // 0x3df8
	13'h1efd: q1 = 16'h610a; // 0x3dfa
	13'h1efe: q1 = 16'h4eb9; // 0x3dfc
	13'h1eff: q1 = 16'h0000; // 0x3dfe
	13'h1f00: q1 = 16'h01d8; // 0x3e00
	13'h1f01: q1 = 16'h4e5e; // 0x3e02
	13'h1f02: q1 = 16'h4e75; // 0x3e04
	13'h1f03: q1 = 16'h4e56; // 0x3e06
	13'h1f04: q1 = 16'hfffe; // 0x3e08
	13'h1f05: q1 = 16'h48e7; // 0x3e0a
	13'h1f06: q1 = 16'h101c; // 0x3e0c
	13'h1f07: q1 = 16'h2a7c; // 0x3e0e
	13'h1f08: q1 = 16'h0001; // 0x3e10
	13'h1f09: q1 = 16'h7b42; // 0x3e12
	13'h1f0a: q1 = 16'h4cf9; // 0x3e14
	13'h1f0b: q1 = 16'h0703; // 0x3e16
	13'h1f0c: q1 = 16'h0001; // 0x3e18
	13'h1f0d: q1 = 16'h77ea; // 0x3e1a
	13'h1f0e: q1 = 16'h48f9; // 0x3e1c
	13'h1f0f: q1 = 16'h0703; // 0x3e1e
	13'h1f10: q1 = 16'h0001; // 0x3e20
	13'h1f11: q1 = 16'h7a1e; // 0x3e22
	13'h1f12: q1 = 16'h4cb9; // 0x3e24
	13'h1f13: q1 = 16'h0703; // 0x3e26
	13'h1f14: q1 = 16'h0001; // 0x3e28
	13'h1f15: q1 = 16'h77fe; // 0x3e2a
	13'h1f16: q1 = 16'h48b9; // 0x3e2c
	13'h1f17: q1 = 16'h0703; // 0x3e2e
	13'h1f18: q1 = 16'h0001; // 0x3e30
	13'h1f19: q1 = 16'h7a32; // 0x3e32
	13'h1f1a: q1 = 16'h206e; // 0x3e34
	13'h1f1b: q1 = 16'h0008; // 0x3e36
	13'h1f1c: q1 = 16'h3d58; // 0x3e38
	13'h1f1d: q1 = 16'hfffe; // 0x3e3a
	13'h1f1e: q1 = 16'h2f08; // 0x3e3c
	13'h1f1f: q1 = 16'h4267; // 0x3e3e
	13'h1f20: q1 = 16'h6100; // 0x3e40
	13'h1f21: q1 = 16'h00dc; // 0x3e42
	13'h1f22: q1 = 16'h4a40; // 0x3e44
	13'h1f23: q1 = 16'h660e; // 0x3e46
	13'h1f24: q1 = 16'h3eae; // 0x3e48
	13'h1f25: q1 = 16'hfffe; // 0x3e4a
	13'h1f26: q1 = 16'h6100; // 0x3e4c
	13'h1f27: q1 = 16'h00d0; // 0x3e4e
	13'h1f28: q1 = 16'h4a40; // 0x3e50
	13'h1f29: q1 = 16'h6700; // 0x3e52
	13'h1f2a: q1 = 16'h00be; // 0x3e54
	13'h1f2b: q1 = 16'h5c8f; // 0x3e56
	13'h1f2c: q1 = 16'h4a90; // 0x3e58
	13'h1f2d: q1 = 16'h6ce0; // 0x3e5a
	13'h1f2e: q1 = 16'h3abc; // 0x3e5c
	13'h1f2f: q1 = 16'hffff; // 0x3e5e
	13'h1f30: q1 = 16'h2a7c; // 0x3e60
	13'h1f31: q1 = 16'h0001; // 0x3e62
	13'h1f32: q1 = 16'h7b42; // 0x3e64
	13'h1f33: q1 = 16'h4a5d; // 0x3e66
	13'h1f34: q1 = 16'h6d00; // 0x3e68
	13'h1f35: q1 = 16'h0090; // 0x3e6a
	13'h1f36: q1 = 16'h361d; // 0x3e6c
	13'h1f37: q1 = 16'h267c; // 0x3e6e
	13'h1f38: q1 = 16'h0001; // 0x3e70
	13'h1f39: q1 = 16'h7a00; // 0x3e72
	13'h1f3a: q1 = 16'h3433; // 0x3e74
	13'h1f3b: q1 = 16'h3000; // 0x3e76
	13'h1f3c: q1 = 16'h6f0a; // 0x3e78
	13'h1f3d: q1 = 16'h3f02; // 0x3e7a
	13'h1f3e: q1 = 16'h4eb9; // 0x3e7c
	13'h1f3f: q1 = 16'h0000; // 0x3e7e
	13'h1f40: q1 = 16'h824a; // 0x3e80
	13'h1f41: q1 = 16'h548f; // 0x3e82
	13'h1f42: q1 = 16'h082d; // 0x3e84
	13'h1f43: q1 = 16'h0000; // 0x3e86
	13'h1f44: q1 = 16'hfffd; // 0x3e88
	13'h1f45: q1 = 16'h674a; // 0x3e8a
	13'h1f46: q1 = 16'h285d; // 0x3e8c
	13'h1f47: q1 = 16'h267c; // 0x3e8e
	13'h1f48: q1 = 16'h0000; // 0x3e90
	13'h1f49: q1 = 16'hca60; // 0x3e92
	13'h1f4a: q1 = 16'h3673; // 0x3e94
	13'h1f4b: q1 = 16'h3000; // 0x3e96
	13'h1f4c: q1 = 16'hd7fc; // 0x3e98
	13'h1f4d: q1 = 16'h0001; // 0x3e9a
	13'h1f4e: q1 = 16'h7808; // 0x3e9c
	13'h1f4f: q1 = 16'h4cd4; // 0x3e9e
	13'h1f50: q1 = 16'h0303; // 0x3ea0
	13'h1f51: q1 = 16'h48d3; // 0x3ea2
	13'h1f52: q1 = 16'h0303; // 0x3ea4
	13'h1f53: q1 = 16'h4cec; // 0x3ea6
	13'h1f54: q1 = 16'h0303; // 0x3ea8
	13'h1f55: q1 = 16'h0010; // 0x3eaa
	13'h1f56: q1 = 16'h48eb; // 0x3eac
	13'h1f57: q1 = 16'h0303; // 0x3eae
	13'h1f58: q1 = 16'h0010; // 0x3eb0
	13'h1f59: q1 = 16'h082d; // 0x3eb2
	13'h1f5a: q1 = 16'h0001; // 0x3eb4
	13'h1f5b: q1 = 16'hfff9; // 0x3eb6
	13'h1f5c: q1 = 16'h6624; // 0x3eb8
	13'h1f5d: q1 = 16'h267c; // 0x3eba
	13'h1f5e: q1 = 16'h0001; // 0x3ebc
	13'h1f5f: q1 = 16'h77ea; // 0x3ebe
	13'h1f60: q1 = 16'h37ae; // 0x3ec0
	13'h1f61: q1 = 16'hfffe; // 0x3ec2
	13'h1f62: q1 = 16'h3000; // 0x3ec4
	13'h1f63: q1 = 16'h267c; // 0x3ec6
	13'h1f64: q1 = 16'h0001; // 0x3ec8
	13'h1f65: q1 = 16'h7a00; // 0x3eca
	13'h1f66: q1 = 16'h37b9; // 0x3ecc
	13'h1f67: q1 = 16'h0001; // 0x3ece
	13'h1f68: q1 = 16'h7a3c; // 0x3ed0
	13'h1f69: q1 = 16'h3000; // 0x3ed2
	13'h1f6a: q1 = 16'h6090; // 0x3ed4
	13'h1f6b: q1 = 16'h082d; // 0x3ed6
	13'h1f6c: q1 = 16'h0001; // 0x3ed8
	13'h1f6d: q1 = 16'hfffd; // 0x3eda
	13'h1f6e: q1 = 16'h67dc; // 0x3edc
	13'h1f6f: q1 = 16'h285d; // 0x3ede
	13'h1f70: q1 = 16'h267c; // 0x3ee0
	13'h1f71: q1 = 16'h0000; // 0x3ee2
	13'h1f72: q1 = 16'hca7e; // 0x3ee4
	13'h1f73: q1 = 16'h3673; // 0x3ee6
	13'h1f74: q1 = 16'h3000; // 0x3ee8
	13'h1f75: q1 = 16'hd7fc; // 0x3eea
	13'h1f76: q1 = 16'h0001; // 0x3eec
	13'h1f77: q1 = 16'h7808; // 0x3eee
	13'h1f78: q1 = 16'h4cd4; // 0x3ef0
	13'h1f79: q1 = 16'h0003; // 0x3ef2
	13'h1f7a: q1 = 16'h48d3; // 0x3ef4
	13'h1f7b: q1 = 16'h0003; // 0x3ef6
	13'h1f7c: q1 = 16'h60c0; // 0x3ef8
	13'h1f7d: q1 = 16'h3039; // 0x3efa
	13'h1f7e: q1 = 16'h0001; // 0x3efc
	13'h1f7f: q1 = 16'h7a3c; // 0x3efe
	13'h1f80: q1 = 16'h5279; // 0x3f00
	13'h1f81: q1 = 16'h0001; // 0x3f02
	13'h1f82: q1 = 16'h7a3c; // 0x3f04
	13'h1f83: q1 = 16'h680e; // 0x3f06
	13'h1f84: q1 = 16'h33fc; // 0x3f08
	13'h1f85: q1 = 16'h0001; // 0x3f0a
	13'h1f86: q1 = 16'h0001; // 0x3f0c
	13'h1f87: q1 = 16'h7a3c; // 0x3f0e
	13'h1f88: q1 = 16'h6004; // 0x3f10
	13'h1f89: q1 = 16'h5c8f; // 0x3f12
	13'h1f8a: q1 = 16'h4240; // 0x3f14
	13'h1f8b: q1 = 16'h4cdf; // 0x3f16
	13'h1f8c: q1 = 16'h3808; // 0x3f18
	13'h1f8d: q1 = 16'h4e5e; // 0x3f1a
	13'h1f8e: q1 = 16'h4e75; // 0x3f1c
	13'h1f8f: q1 = 16'h4e56; // 0x3f1e
	13'h1f90: q1 = 16'h0000; // 0x3f20
	13'h1f91: q1 = 16'h206e; // 0x3f22
	13'h1f92: q1 = 16'h000a; // 0x3f24
	13'h1f93: q1 = 16'h3018; // 0x3f26
	13'h1f94: q1 = 16'he540; // 0x3f28
	13'h1f95: q1 = 16'h247c; // 0x3f2a
	13'h1f96: q1 = 16'h0000; // 0x3f2c
	13'h1f97: q1 = 16'hf4f6; // 0x3f2e
	13'h1f98: q1 = 16'h2472; // 0x3f30
	13'h1f99: q1 = 16'h0000; // 0x3f32
	13'h1f9a: q1 = 16'h4e92; // 0x3f34
	13'h1f9b: q1 = 16'h4e5e; // 0x3f36
	13'h1f9c: q1 = 16'h4e75; // 0x3f38
	13'h1f9d: q1 = 16'h247c; // 0x3f3a
	13'h1f9e: q1 = 16'h0000; // 0x3f3c
	13'h1f9f: q1 = 16'hf506; // 0x3f3e
	13'h1fa0: q1 = 16'h6100; // 0x3f40
	13'h1fa1: q1 = 16'h006c; // 0x3f42
	13'h1fa2: q1 = 16'h4a40; // 0x3f44
	13'h1fa3: q1 = 16'h6602; // 0x3f46
	13'h1fa4: q1 = 16'h4e75; // 0x3f48
	13'h1fa5: q1 = 16'h6100; // 0x3f4a
	13'h1fa6: q1 = 16'h0080; // 0x3f4c
	13'h1fa7: q1 = 16'h3afc; // 0x3f4e
	13'h1fa8: q1 = 16'h0001; // 0x3f50
	13'h1fa9: q1 = 16'h3ac2; // 0x3f52
	13'h1faa: q1 = 16'h2ad8; // 0x3f54
	13'h1fab: q1 = 16'h7001; // 0x3f56
	13'h1fac: q1 = 16'h4e75; // 0x3f58
	13'h1fad: q1 = 16'h247c; // 0x3f5a
	13'h1fae: q1 = 16'h0000; // 0x3f5c
	13'h1faf: q1 = 16'hf514; // 0x3f5e
	13'h1fb0: q1 = 16'h614c; // 0x3f60
	13'h1fb1: q1 = 16'h4a40; // 0x3f62
	13'h1fb2: q1 = 16'h6602; // 0x3f64
	13'h1fb3: q1 = 16'h4e75; // 0x3f66
	13'h1fb4: q1 = 16'h6162; // 0x3f68
	13'h1fb5: q1 = 16'h3afc; // 0x3f6a
	13'h1fb6: q1 = 16'h0003; // 0x3f6c
	13'h1fb7: q1 = 16'h3ac2; // 0x3f6e
	13'h1fb8: q1 = 16'h2ad8; // 0x3f70
	13'h1fb9: q1 = 16'h2ad8; // 0x3f72
	13'h1fba: q1 = 16'h7001; // 0x3f74
	13'h1fbb: q1 = 16'h4e75; // 0x3f76
	13'h1fbc: q1 = 16'h4e75; // 0x3f78
	13'h1fbd: q1 = 16'h247c; // 0x3f7a
	13'h1fbe: q1 = 16'h0000; // 0x3f7c
	13'h1fbf: q1 = 16'hf514; // 0x3f7e
	13'h1fc0: q1 = 16'h612c; // 0x3f80
	13'h1fc1: q1 = 16'h4a40; // 0x3f82
	13'h1fc2: q1 = 16'h6726; // 0x3f84
	13'h1fc3: q1 = 16'h3231; // 0x3f86
	13'h1fc4: q1 = 16'h2002; // 0x3f88
	13'h1fc5: q1 = 16'h4a41; // 0x3f8a
	13'h1fc6: q1 = 16'h670a; // 0x3f8c
	13'h1fc7: q1 = 16'hb26e; // 0x3f8e
	13'h1fc8: q1 = 16'h0008; // 0x3f90
	13'h1fc9: q1 = 16'h6d04; // 0x3f92
	13'h1fca: q1 = 16'h611e; // 0x3f94
	13'h1fcb: q1 = 16'h60ea; // 0x3f96
	13'h1fcc: q1 = 16'h2258; // 0x3f98
	13'h1fcd: q1 = 16'h3282; // 0x3f9a
	13'h1fce: q1 = 16'h425d; // 0x3f9c
	13'h1fcf: q1 = 16'h3ac2; // 0x3f9e
	13'h1fd0: q1 = 16'h612a; // 0x3fa0
	13'h1fd1: q1 = 16'h5442; // 0x3fa2
	13'h1fd2: q1 = 16'h425d; // 0x3fa4
	13'h1fd3: q1 = 16'h3ac2; // 0x3fa6
	13'h1fd4: q1 = 16'h6122; // 0x3fa8
	13'h1fd5: q1 = 16'h7001; // 0x3faa
	13'h1fd6: q1 = 16'h4e75; // 0x3fac
	13'h1fd7: q1 = 16'h227c; // 0x3fae
	13'h1fd8: q1 = 16'h0001; // 0x3fb0
	13'h1fd9: q1 = 16'h7a1e; // 0x3fb2
	13'h1fda: q1 = 16'h141a; // 0x3fb4
	13'h1fdb: q1 = 16'h6d10; // 0x3fb6
	13'h1fdc: q1 = 16'h4882; // 0x3fb8
	13'h1fdd: q1 = 16'h3231; // 0x3fba
	13'h1fde: q1 = 16'h2000; // 0x3fbc
	13'h1fdf: q1 = 16'hb26e; // 0x3fbe
	13'h1fe0: q1 = 16'h0008; // 0x3fc0
	13'h1fe1: q1 = 16'h6ef0; // 0x3fc2
	13'h1fe2: q1 = 16'h7001; // 0x3fc4
	13'h1fe3: q1 = 16'h4e75; // 0x3fc6
	13'h1fe4: q1 = 16'h4240; // 0x3fc8
	13'h1fe5: q1 = 16'h4e75; // 0x3fca
	13'h1fe6: q1 = 16'h247c; // 0x3fcc
	13'h1fe7: q1 = 16'h0001; // 0x3fce
	13'h1fe8: q1 = 16'h7a00; // 0x3fd0
	13'h1fe9: q1 = 16'h3032; // 0x3fd2
	13'h1fea: q1 = 16'h2000; // 0x3fd4
	13'h1feb: q1 = 16'h6718; // 0x3fd6
	13'h1fec: q1 = 16'h721c; // 0x3fd8
	13'h1fed: q1 = 16'hb072; // 0x3fda
	13'h1fee: q1 = 16'h1000; // 0x3fdc
	13'h1fef: q1 = 16'h660c; // 0x3fde
	13'h1ff0: q1 = 16'h0c72; // 0x3fe0
	13'h1ff1: q1 = 16'h7fff; // 0x3fe2
	13'h1ff2: q1 = 16'h101e; // 0x3fe4
	13'h1ff3: q1 = 16'h6708; // 0x3fe6
	13'h1ff4: q1 = 16'h4272; // 0x3fe8
	13'h1ff5: q1 = 16'h101e; // 0x3fea
	13'h1ff6: q1 = 16'h5541; // 0x3fec
	13'h1ff7: q1 = 16'h6cea; // 0x3fee
	13'h1ff8: q1 = 16'h35bc; // 0x3ff0
	13'h1ff9: q1 = 16'h7fff; // 0x3ff2
	13'h1ffa: q1 = 16'h201e; // 0x3ff4
	13'h1ffb: q1 = 16'h4e75; // 0x3ff6
	13'h1ffc: q1 = 16'h3039; // 0x3ff8
	13'h1ffd: q1 = 16'h0001; // 0x3ffa
	13'h1ffe: q1 = 16'h7fc6; // 0x3ffc
	13'h1fff: q1 = 16'h6704; // 0x3ffe
  endcase

  always @(posedge clk)
    case (a)
	// foodfight code 136020-306.9e, 136020-305.8e
	13'h0000: q2 = 16'h4240; // 0x0000
	13'h0001: q2 = 16'h4e75; // 0x0002
	13'h0002: q2 = 16'h4e56; // 0x0004
	13'h0003: q2 = 16'h0000; // 0x0006
	13'h0004: q2 = 16'h207c; // 0x0008
	13'h0005: q2 = 16'h0001; // 0x000a
	13'h0006: q2 = 16'h7a3e; // 0x000c
	13'h0007: q2 = 16'h4aa8; // 0x000e
	13'h0008: q2 = 16'h000e; // 0x0010
	13'h0009: q2 = 16'h6710; // 0x0012
	13'h000a: q2 = 16'hd0fc; // 0x0014
	13'h000b: q2 = 16'h0082; // 0x0016
	13'h000c: q2 = 16'h4aa8; // 0x0018
	13'h000d: q2 = 16'h000e; // 0x001a
	13'h000e: q2 = 16'h6706; // 0x001c
	13'h000f: q2 = 16'h4240; // 0x001e
	13'h0010: q2 = 16'h4e5e; // 0x0020
	13'h0011: q2 = 16'h4e75; // 0x0022
	13'h0012: q2 = 16'h42a8; // 0x0024
	13'h0013: q2 = 16'h0000; // 0x0026
	13'h0014: q2 = 16'h4268; // 0x0028
	13'h0015: q2 = 16'h0004; // 0x002a
	13'h0016: q2 = 16'h42a8; // 0x002c
	13'h0017: q2 = 16'h0006; // 0x002e
	13'h0018: q2 = 16'h42a8; // 0x0030
	13'h0019: q2 = 16'h000a; // 0x0032
	13'h001a: q2 = 16'h217c; // 0x0034
	13'h001b: q2 = 16'h0000; // 0x0036
	13'h001c: q2 = 16'hbba4; // 0x0038
	13'h001d: q2 = 16'h0012; // 0x003a
	13'h001e: q2 = 16'h216e; // 0x003c
	13'h001f: q2 = 16'h0008; // 0x003e
	13'h0020: q2 = 16'h000e; // 0x0040
	13'h0021: q2 = 16'h2008; // 0x0042
	13'h0022: q2 = 16'h4e5e; // 0x0044
	13'h0023: q2 = 16'h4e75; // 0x0046
	13'h0024: q2 = 16'h5279; // 0x0048
	13'h0025: q2 = 16'h0001; // 0x004a
	13'h0026: q2 = 16'h7b9c; // 0x004c
	13'h0027: q2 = 16'h6706; // 0x004e
	13'h0028: q2 = 16'h4e71; // 0x0050
	13'h0029: q2 = 16'h4e71; // 0x0052
	13'h002a: q2 = 16'h4e75; // 0x0054
	13'h002b: q2 = 16'h48e7; // 0x0056
	13'h002c: q2 = 16'h0610; // 0x0058
	13'h002d: q2 = 16'h2479; // 0x005a
	13'h002e: q2 = 16'h0000; // 0x005c
	13'h002f: q2 = 16'hf51c; // 0x005e
	13'h0030: q2 = 16'h267c; // 0x0060
	13'h0031: q2 = 16'h0001; // 0x0062
	13'h0032: q2 = 16'h7808; // 0x0064
	13'h0033: q2 = 16'h4245; // 0x0066
	13'h0034: q2 = 16'h7c03; // 0x0068
	13'h0035: q2 = 16'h2013; // 0x006a
	13'h0036: q2 = 16'h2040; // 0x006c
	13'h0037: q2 = 16'h6706; // 0x006e
	13'h0038: q2 = 16'h4e90; // 0x0070
	13'h0039: q2 = 16'hee40; // 0x0072
	13'h003a: q2 = 16'h3480; // 0x0074
	13'h003b: q2 = 16'h548a; // 0x0076
	13'h003c: q2 = 16'hd7fc; // 0x0078
	13'h003d: q2 = 16'h0000; // 0x007a
	13'h003e: q2 = 16'h000c; // 0x007c
	13'h003f: q2 = 16'h2013; // 0x007e
	13'h0040: q2 = 16'h2040; // 0x0080
	13'h0041: q2 = 16'h6700; // 0x0082
	13'h0042: q2 = 16'h00a8; // 0x0084
	13'h0043: q2 = 16'h4e90; // 0x0086
	13'h0044: q2 = 16'h6608; // 0x0088
	13'h0045: q2 = 16'h6100; // 0x008a
	13'h0046: q2 = 16'h0146; // 0x008c
	13'h0047: q2 = 16'h6000; // 0x008e
	13'h0048: q2 = 16'h009c; // 0x0090
	13'h0049: q2 = 16'hee48; // 0x0092
	13'h004a: q2 = 16'hd7fc; // 0x0094
	13'h004b: q2 = 16'h0000; // 0x0096
	13'h004c: q2 = 16'h000c; // 0x0098
	13'h004d: q2 = 16'h2413; // 0x009a
	13'h004e: q2 = 16'h2042; // 0x009c
	13'h004f: q2 = 16'h6700; // 0x009e
	13'h0050: q2 = 16'h0084; // 0x00a0
	13'h0051: q2 = 16'h6100; // 0x00a2
	13'h0052: q2 = 16'h0108; // 0x00a4
	13'h0053: q2 = 16'h3480; // 0x00a6
	13'h0054: q2 = 16'h508b; // 0x00a8
	13'h0055: q2 = 16'h548a; // 0x00aa
	13'h0056: q2 = 16'h51ce; // 0x00ac
	13'h0057: q2 = 16'hffbc; // 0x00ae
	13'h0058: q2 = 16'h4240; // 0x00b0
	13'h0059: q2 = 16'h2213; // 0x00b2
	13'h005a: q2 = 16'h2041; // 0x00b4
	13'h005b: q2 = 16'h6704; // 0x00b6
	13'h005c: q2 = 16'h6100; // 0x00b8
	13'h005d: q2 = 16'h00f2; // 0x00ba
	13'h005e: q2 = 16'he348; // 0x00bc
	13'h005f: q2 = 16'h508b; // 0x00be
	13'h0060: q2 = 16'h2213; // 0x00c0
	13'h0061: q2 = 16'h2041; // 0x00c2
	13'h0062: q2 = 16'h6704; // 0x00c4
	13'h0063: q2 = 16'h6100; // 0x00c6
	13'h0064: q2 = 16'h00e4; // 0x00c8
	13'h0065: q2 = 16'h508b; // 0x00ca
	13'h0066: q2 = 16'h2213; // 0x00cc
	13'h0067: q2 = 16'h2041; // 0x00ce
	13'h0068: q2 = 16'h6704; // 0x00d0
	13'h0069: q2 = 16'h6100; // 0x00d2
	13'h006a: q2 = 16'h00d8; // 0x00d4
	13'h006b: q2 = 16'he348; // 0x00d6
	13'h006c: q2 = 16'h508b; // 0x00d8
	13'h006d: q2 = 16'h2213; // 0x00da
	13'h006e: q2 = 16'h2041; // 0x00dc
	13'h006f: q2 = 16'h6704; // 0x00de
	13'h0070: q2 = 16'h6100; // 0x00e0
	13'h0071: q2 = 16'h00ca; // 0x00e2
	13'h0072: q2 = 16'he448; // 0x00e4
	13'h0073: q2 = 16'h508b; // 0x00e6
	13'h0074: q2 = 16'h2213; // 0x00e8
	13'h0075: q2 = 16'h2041; // 0x00ea
	13'h0076: q2 = 16'h6710; // 0x00ec
	13'h0077: q2 = 16'h6100; // 0x00ee
	13'h0078: q2 = 16'h00bc; // 0x00f0
	13'h0079: q2 = 16'h660a; // 0x00f2
	13'h007a: q2 = 16'h3400; // 0x00f4
	13'h007b: q2 = 16'h6100; // 0x00f6
	13'h007c: q2 = 16'h00da; // 0x00f8
	13'h007d: q2 = 16'h3002; // 0x00fa
	13'h007e: q2 = 16'h6002; // 0x00fc
	13'h007f: q2 = 16'h3480; // 0x00fe
	13'h0080: q2 = 16'hba7c; // 0x0100
	13'h0081: q2 = 16'h0014; // 0x0102
	13'h0082: q2 = 16'h6714; // 0x0104
	13'h0083: q2 = 16'h508b; // 0x0106
	13'h0084: q2 = 16'h94fc; // 0x0108
	13'h0085: q2 = 16'h0010; // 0x010a
	13'h0086: q2 = 16'hd5f9; // 0x010c
	13'h0087: q2 = 16'h0000; // 0x010e
	13'h0088: q2 = 16'hf520; // 0x0110
	13'h0089: q2 = 16'hda7c; // 0x0112
	13'h008a: q2 = 16'h000a; // 0x0114
	13'h008b: q2 = 16'h6000; // 0x0116
	13'h008c: q2 = 16'hff50; // 0x0118
	13'h008d: q2 = 16'h4cdf; // 0x011a
	13'h008e: q2 = 16'h0860; // 0x011c
	13'h008f: q2 = 16'h4ef9; // 0x011e
	13'h0090: q2 = 16'h0000; // 0x0120
	13'h0091: q2 = 16'hba38; // 0x0122
	13'h0092: q2 = 16'h807c; // 0x0124
	13'h0093: q2 = 16'h00e0; // 0x0126
	13'h0094: q2 = 16'h6000; // 0x0128
	13'h0095: q2 = 16'hff7c; // 0x012a
	13'h0096: q2 = 16'hd7fc; // 0x012c
	13'h0097: q2 = 16'h0000; // 0x012e
	13'h0098: q2 = 16'h0014; // 0x0130
	13'h0099: q2 = 16'h6000; // 0x0132
	13'h009a: q2 = 16'hff76; // 0x0134
	13'h009b: q2 = 16'h4a6b; // 0x0136
	13'h009c: q2 = 16'h000a; // 0x0138
	13'h009d: q2 = 16'h6606; // 0x013a
	13'h009e: q2 = 16'h26bc; // 0x013c
	13'h009f: q2 = 16'h0000; // 0x013e
	13'h00a0: q2 = 16'h8150; // 0x0140
	13'h00a1: q2 = 16'h536b; // 0x0142
	13'h00a2: q2 = 16'h000a; // 0x0144
	13'h00a3: q2 = 16'h302b; // 0x0146
	13'h00a4: q2 = 16'h0008; // 0x0148
	13'h00a5: q2 = 16'h44fc; // 0x014a
	13'h00a6: q2 = 16'h0000; // 0x014c
	13'h00a7: q2 = 16'h4e75; // 0x014e
	13'h00a8: q2 = 16'h206b; // 0x0150
	13'h00a9: q2 = 16'h0004; // 0x0152
	13'h00aa: q2 = 16'h3768; // 0x0154
	13'h00ab: q2 = 16'h0004; // 0x0156
	13'h00ac: q2 = 16'h000a; // 0x0158
	13'h00ad: q2 = 16'h6e16; // 0x015a
	13'h00ae: q2 = 16'h670c; // 0x015c
	13'h00af: q2 = 16'h302b; // 0x015e
	13'h00b0: q2 = 16'h000a; // 0x0160
	13'h00b1: q2 = 16'h48c0; // 0x0162
	13'h00b2: q2 = 16'hd1ab; // 0x0164
	13'h00b3: q2 = 16'h0004; // 0x0166
	13'h00b4: q2 = 16'h60e6; // 0x0168
	13'h00b5: q2 = 16'h302b; // 0x016a
	13'h00b6: q2 = 16'h0008; // 0x016c
	13'h00b7: q2 = 16'h4293; // 0x016e
	13'h00b8: q2 = 16'h4e75; // 0x0170
	13'h00b9: q2 = 16'h3010; // 0x0172
	13'h00ba: q2 = 16'hd06b; // 0x0174
	13'h00bb: q2 = 16'h0008; // 0x0176
	13'h00bc: q2 = 16'h3740; // 0x0178
	13'h00bd: q2 = 16'h0008; // 0x017a
	13'h00be: q2 = 16'h54ab; // 0x017c
	13'h00bf: q2 = 16'h0004; // 0x017e
	13'h00c0: q2 = 16'h26bc; // 0x0180
	13'h00c1: q2 = 16'h0000; // 0x0182
	13'h00c2: q2 = 16'h819c; // 0x0184
	13'h00c3: q2 = 16'h536b; // 0x0186
	13'h00c4: q2 = 16'h000a; // 0x0188
	13'h00c5: q2 = 16'h660e; // 0x018a
	13'h00c6: q2 = 16'h58ab; // 0x018c
	13'h00c7: q2 = 16'h0004; // 0x018e
	13'h00c8: q2 = 16'h26bc; // 0x0190
	13'h00c9: q2 = 16'h0000; // 0x0192
	13'h00ca: q2 = 16'h8150; // 0x0194
	13'h00cb: q2 = 16'h44fc; // 0x0196
	13'h00cc: q2 = 16'h0000; // 0x0198
	13'h00cd: q2 = 16'h4e75; // 0x019a
	13'h00ce: q2 = 16'h206b; // 0x019c
	13'h00cf: q2 = 16'h0004; // 0x019e
	13'h00d0: q2 = 16'h3010; // 0x01a0
	13'h00d1: q2 = 16'hd06b; // 0x01a2
	13'h00d2: q2 = 16'h0008; // 0x01a4
	13'h00d3: q2 = 16'h3740; // 0x01a6
	13'h00d4: q2 = 16'h0008; // 0x01a8
	13'h00d5: q2 = 16'h60da; // 0x01aa
	13'h00d6: q2 = 16'h4a6b; // 0x01ac
	13'h00d7: q2 = 16'h0006; // 0x01ae
	13'h00d8: q2 = 16'h6612; // 0x01b0
	13'h00d9: q2 = 16'h2253; // 0x01b2
	13'h00da: q2 = 16'h3759; // 0x01b4
	13'h00db: q2 = 16'h0004; // 0x01b6
	13'h00dc: q2 = 16'h3759; // 0x01b8
	13'h00dd: q2 = 16'h0006; // 0x01ba
	13'h00de: q2 = 16'h6604; // 0x01bc
	13'h00df: q2 = 16'h4293; // 0x01be
	13'h00e0: q2 = 16'h4e75; // 0x01c0
	13'h00e1: q2 = 16'h2689; // 0x01c2
	13'h00e2: q2 = 16'h806b; // 0x01c4
	13'h00e3: q2 = 16'h0004; // 0x01c6
	13'h00e4: q2 = 16'h536b; // 0x01c8
	13'h00e5: q2 = 16'h0006; // 0x01ca
	13'h00e6: q2 = 16'h44fc; // 0x01cc
	13'h00e7: q2 = 16'h0000; // 0x01ce
	13'h00e8: q2 = 16'h4e75; // 0x01d0
	13'h00e9: q2 = 16'h300a; // 0x01d2
	13'h00ea: q2 = 16'he248; // 0x01d4
	13'h00eb: q2 = 16'hc07c; // 0x01d6
	13'h00ec: q2 = 16'h000e; // 0x01d8
	13'h00ed: q2 = 16'hd045; // 0x01da
	13'h00ee: q2 = 16'h6102; // 0x01dc
	13'h00ef: q2 = 16'h4e75; // 0x01de
	13'h00f0: q2 = 16'h227c; // 0x01e0
	13'h00f1: q2 = 16'h0000; // 0x01e2
	13'h00f2: q2 = 16'hca60; // 0x01e4
	13'h00f3: q2 = 16'hd2c0; // 0x01e6
	13'h00f4: q2 = 16'h3211; // 0x01e8
	13'h00f5: q2 = 16'h6d36; // 0x01ea
	13'h00f6: q2 = 16'h227c; // 0x01ec
	13'h00f7: q2 = 16'h0001; // 0x01ee
	13'h00f8: q2 = 16'h7808; // 0x01f0
	13'h00f9: q2 = 16'hd2c1; // 0x01f2
	13'h00fa: q2 = 16'h4291; // 0x01f4
	13'h00fb: q2 = 16'h42a9; // 0x01f6
	13'h00fc: q2 = 16'h000c; // 0x01f8
	13'h00fd: q2 = 16'h42a9; // 0x01fa
	13'h00fe: q2 = 16'h0018; // 0x01fc
	13'h00ff: q2 = 16'h3200; // 0x01fe
	13'h0100: q2 = 16'h2279; // 0x0200
	13'h0101: q2 = 16'h0000; // 0x0202
	13'h0102: q2 = 16'hf51c; // 0x0204
	13'h0103: q2 = 16'h5449; // 0x0206
	13'h0104: q2 = 16'hb27c; // 0x0208
	13'h0105: q2 = 16'h000a; // 0x020a
	13'h0106: q2 = 16'h6d0c; // 0x020c
	13'h0107: q2 = 16'hd3f9; // 0x020e
	13'h0108: q2 = 16'h0000; // 0x0210
	13'h0109: q2 = 16'hf520; // 0x0212
	13'h010a: q2 = 16'h927c; // 0x0214
	13'h010b: q2 = 16'h000a; // 0x0216
	13'h010c: q2 = 16'h60ee; // 0x0218
	13'h010d: q2 = 16'he349; // 0x021a
	13'h010e: q2 = 16'h33bc; // 0x021c
	13'h010f: q2 = 16'h00e0; // 0x021e
	13'h0110: q2 = 16'h1000; // 0x0220
	13'h0111: q2 = 16'h227c; // 0x0222
	13'h0112: q2 = 16'h0000; // 0x0224
	13'h0113: q2 = 16'hca7e; // 0x0226
	13'h0114: q2 = 16'hd2c0; // 0x0228
	13'h0115: q2 = 16'h3251; // 0x022a
	13'h0116: q2 = 16'hd3fc; // 0x022c
	13'h0117: q2 = 16'h0001; // 0x022e
	13'h0118: q2 = 16'h7808; // 0x0230
	13'h0119: q2 = 16'h4291; // 0x0232
	13'h011a: q2 = 16'h227c; // 0x0234
	13'h011b: q2 = 16'h0001; // 0x0236
	13'h011c: q2 = 16'h7a00; // 0x0238
	13'h011d: q2 = 16'hd2c0; // 0x023a
	13'h011e: q2 = 16'h4251; // 0x023c
	13'h011f: q2 = 16'h227c; // 0x023e
	13'h0120: q2 = 16'h0001; // 0x0240
	13'h0121: q2 = 16'h77ea; // 0x0242
	13'h0122: q2 = 16'hd2c0; // 0x0244
	13'h0123: q2 = 16'h4251; // 0x0246
	13'h0124: q2 = 16'h4e75; // 0x0248
	13'h0125: q2 = 16'h4e56; // 0x024a
	13'h0126: q2 = 16'h0000; // 0x024c
	13'h0127: q2 = 16'h2f03; // 0x024e
	13'h0128: q2 = 16'h362e; // 0x0250
	13'h0129: q2 = 16'h0008; // 0x0252
	13'h012a: q2 = 16'h701c; // 0x0254
	13'h012b: q2 = 16'h207c; // 0x0256
	13'h012c: q2 = 16'h0001; // 0x0258
	13'h012d: q2 = 16'h7a00; // 0x025a
	13'h012e: q2 = 16'hb670; // 0x025c
	13'h012f: q2 = 16'h0000; // 0x025e
	13'h0130: q2 = 16'h6606; // 0x0260
	13'h0131: q2 = 16'h4e71; // 0x0262
	13'h0132: q2 = 16'h6100; // 0x0264
	13'h0133: q2 = 16'hff7a; // 0x0266
	13'h0134: q2 = 16'h4a40; // 0x0268
	13'h0135: q2 = 16'h6704; // 0x026a
	13'h0136: q2 = 16'h5540; // 0x026c
	13'h0137: q2 = 16'h60ec; // 0x026e
	13'h0138: q2 = 16'h261f; // 0x0270
	13'h0139: q2 = 16'h4e5e; // 0x0272
	13'h013a: q2 = 16'h4e75; // 0x0274
	13'h013b: q2 = 16'h5693; // 0x0276
	13'h013c: q2 = 16'hdc24; // 0x0278
	13'h013d: q2 = 16'h6bd5; // 0x027a
	13'h013e: q2 = 16'h7398; // 0x027c
	13'h013f: q2 = 16'h4e56; // 0x027e
	13'h0140: q2 = 16'hfffc; // 0x0280
	13'h0141: q2 = 16'h0c79; // 0x0282
	13'h0142: q2 = 16'h0001; // 0x0284
	13'h0143: q2 = 16'h0001; // 0x0286
	13'h0144: q2 = 16'h87dc; // 0x0288
	13'h0145: q2 = 16'h660a; // 0x028a
	13'h0146: q2 = 16'h4257; // 0x028c
	13'h0147: q2 = 16'h4eb9; // 0x028e
	13'h0148: q2 = 16'h0000; // 0x0290
	13'h0149: q2 = 16'hbdaa; // 0x0292
	13'h014a: q2 = 16'h6034; // 0x0294
	13'h014b: q2 = 16'h2039; // 0x0296
	13'h014c: q2 = 16'h0001; // 0x0298
	13'h014d: q2 = 16'h862c; // 0x029a
	13'h014e: q2 = 16'hb0b9; // 0x029c
	13'h014f: q2 = 16'h0001; // 0x029e
	13'h0150: q2 = 16'h8652; // 0x02a0
	13'h0151: q2 = 16'h6f14; // 0x02a2
	13'h0152: q2 = 16'h4257; // 0x02a4
	13'h0153: q2 = 16'h4eb9; // 0x02a6
	13'h0154: q2 = 16'h0000; // 0x02a8
	13'h0155: q2 = 16'hbdaa; // 0x02aa
	13'h0156: q2 = 16'h3ebc; // 0x02ac
	13'h0157: q2 = 16'h0001; // 0x02ae
	13'h0158: q2 = 16'h4eb9; // 0x02b0
	13'h0159: q2 = 16'h0000; // 0x02b2
	13'h015a: q2 = 16'hbdaa; // 0x02b4
	13'h015b: q2 = 16'h6012; // 0x02b6
	13'h015c: q2 = 16'h3ebc; // 0x02b8
	13'h015d: q2 = 16'h0001; // 0x02ba
	13'h015e: q2 = 16'h4eb9; // 0x02bc
	13'h015f: q2 = 16'h0000; // 0x02be
	13'h0160: q2 = 16'hbdaa; // 0x02c0
	13'h0161: q2 = 16'h4257; // 0x02c2
	13'h0162: q2 = 16'h4eb9; // 0x02c4
	13'h0163: q2 = 16'h0000; // 0x02c6
	13'h0164: q2 = 16'hbdaa; // 0x02c8
	13'h0165: q2 = 16'h4e5e; // 0x02ca
	13'h0166: q2 = 16'h4e75; // 0x02cc
	13'h0167: q2 = 16'h4e56; // 0x02ce
	13'h0168: q2 = 16'h0000; // 0x02d0
	13'h0169: q2 = 16'h48e7; // 0x02d2
	13'h016a: q2 = 16'h0f04; // 0x02d4
	13'h016b: q2 = 16'h3e2e; // 0x02d6
	13'h016c: q2 = 16'h0008; // 0x02d8
	13'h016d: q2 = 16'h3c2e; // 0x02da
	13'h016e: q2 = 16'h000a; // 0x02dc
	13'h016f: q2 = 16'h4257; // 0x02de
	13'h0170: q2 = 16'h3f06; // 0x02e0
	13'h0171: q2 = 16'h3f07; // 0x02e2
	13'h0172: q2 = 16'h4eb9; // 0x02e4
	13'h0173: q2 = 16'h0000; // 0x02e6
	13'h0174: q2 = 16'h8744; // 0x02e8
	13'h0175: q2 = 16'h4a9f; // 0x02ea
	13'h0176: q2 = 16'h3a00; // 0x02ec
	13'h0177: q2 = 16'h4a45; // 0x02ee
	13'h0178: q2 = 16'h6604; // 0x02f0
	13'h0179: q2 = 16'h4240; // 0x02f2
	13'h017a: q2 = 16'h6030; // 0x02f4
	13'h017b: q2 = 16'h3005; // 0x02f6
	13'h017c: q2 = 16'h5340; // 0x02f8
	13'h017d: q2 = 16'he940; // 0x02fa
	13'h017e: q2 = 16'h48c0; // 0x02fc
	13'h017f: q2 = 16'h2a40; // 0x02fe
	13'h0180: q2 = 16'hdbfc; // 0x0300
	13'h0181: q2 = 16'h0001; // 0x0302
	13'h0182: q2 = 16'h893e; // 0x0304
	13'h0183: q2 = 16'h0c6d; // 0x0306
	13'h0184: q2 = 16'h0005; // 0x0308
	13'h0185: q2 = 16'h0004; // 0x030a
	13'h0186: q2 = 16'h6714; // 0x030c
	13'h0187: q2 = 16'h536d; // 0x030e
	13'h0188: q2 = 16'h0006; // 0x0310
	13'h0189: q2 = 16'h2e8d; // 0x0312
	13'h018a: q2 = 16'h4eb9; // 0x0314
	13'h018b: q2 = 16'h0000; // 0x0316
	13'h018c: q2 = 16'h161a; // 0x0318
	13'h018d: q2 = 16'h2e8d; // 0x031a
	13'h018e: q2 = 16'h4eb9; // 0x031c
	13'h018f: q2 = 16'h0000; // 0x031e
	13'h0190: q2 = 16'h0f60; // 0x0320
	13'h0191: q2 = 16'h302d; // 0x0322
	13'h0192: q2 = 16'h0004; // 0x0324
	13'h0193: q2 = 16'h4a9f; // 0x0326
	13'h0194: q2 = 16'h4cdf; // 0x0328
	13'h0195: q2 = 16'h20e0; // 0x032a
	13'h0196: q2 = 16'h4e5e; // 0x032c
	13'h0197: q2 = 16'h4e75; // 0x032e
	13'h0198: q2 = 16'h4e56; // 0x0330
	13'h0199: q2 = 16'hfffa; // 0x0332
	13'h019a: q2 = 16'h48e7; // 0x0334
	13'h019b: q2 = 16'h0f0c; // 0x0336
	13'h019c: q2 = 16'h2879; // 0x0338
	13'h019d: q2 = 16'h0001; // 0x033a
	13'h019e: q2 = 16'h7fb8; // 0x033c
	13'h019f: q2 = 16'h2a7c; // 0x033e
	13'h01a0: q2 = 16'h0001; // 0x0340
	13'h01a1: q2 = 16'h893e; // 0x0342
	13'h01a2: q2 = 16'h4247; // 0x0344
	13'h01a3: q2 = 16'hbe7c; // 0x0346
	13'h01a4: q2 = 16'h0008; // 0x0348
	13'h01a5: q2 = 16'h6c10; // 0x034a
	13'h01a6: q2 = 16'h4255; // 0x034c
	13'h01a7: q2 = 16'h426d; // 0x034e
	13'h01a8: q2 = 16'h0002; // 0x0350
	13'h01a9: q2 = 16'hdbfc; // 0x0352
	13'h01aa: q2 = 16'h0000; // 0x0354
	13'h01ab: q2 = 16'h0010; // 0x0356
	13'h01ac: q2 = 16'h5247; // 0x0358
	13'h01ad: q2 = 16'h60ea; // 0x035a
	13'h01ae: q2 = 16'h3014; // 0x035c
	13'h01af: q2 = 16'h5440; // 0x035e
	13'h01b0: q2 = 16'h33c0; // 0x0360
	13'h01b1: q2 = 16'h0001; // 0x0362
	13'h01b2: q2 = 16'h7fa8; // 0x0364
	13'h01b3: q2 = 16'h0c79; // 0x0366
	13'h01b4: q2 = 16'h0008; // 0x0368
	13'h01b5: q2 = 16'h0001; // 0x036a
	13'h01b6: q2 = 16'h7fa8; // 0x036c
	13'h01b7: q2 = 16'h6f08; // 0x036e
	13'h01b8: q2 = 16'h33fc; // 0x0370
	13'h01b9: q2 = 16'h0008; // 0x0372
	13'h01ba: q2 = 16'h0001; // 0x0374
	13'h01bb: q2 = 16'h7fa8; // 0x0376
	13'h01bc: q2 = 16'h3039; // 0x0378
	13'h01bd: q2 = 16'h0001; // 0x037a
	13'h01be: q2 = 16'h7fa8; // 0x037c
	13'h01bf: q2 = 16'hc1fc; // 0x037e
	13'h01c0: q2 = 16'h0005; // 0x0380
	13'h01c1: q2 = 16'h3a00; // 0x0382
	13'h01c2: q2 = 16'h0c54; // 0x0384
	13'h01c3: q2 = 16'h007d; // 0x0386
	13'h01c4: q2 = 16'h6642; // 0x0388
	13'h01c5: q2 = 16'h4a6c; // 0x038a
	13'h01c6: q2 = 16'h0024; // 0x038c
	13'h01c7: q2 = 16'h6c1e; // 0x038e
	13'h01c8: q2 = 16'h3ebc; // 0x0390
	13'h01c9: q2 = 16'h0009; // 0x0392
	13'h01ca: q2 = 16'h4267; // 0x0394
	13'h01cb: q2 = 16'h4eb9; // 0x0396
	13'h01cc: q2 = 16'h0000; // 0x0398
	13'h01cd: q2 = 16'h8e6c; // 0x039a
	13'h01ce: q2 = 16'h4a5f; // 0x039c
	13'h01cf: q2 = 16'h33c0; // 0x039e
	13'h01d0: q2 = 16'h0001; // 0x03a0
	13'h01d1: q2 = 16'h8070; // 0x03a2
	13'h01d2: q2 = 16'h3979; // 0x03a4
	13'h01d3: q2 = 16'h0001; // 0x03a6
	13'h01d4: q2 = 16'h8070; // 0x03a8
	13'h01d5: q2 = 16'h0024; // 0x03aa
	13'h01d6: q2 = 16'h601c; // 0x03ac
	13'h01d7: q2 = 16'h3ebc; // 0x03ae
	13'h01d8: q2 = 16'h0009; // 0x03b0
	13'h01d9: q2 = 16'h4267; // 0x03b2
	13'h01da: q2 = 16'h4eb9; // 0x03b4
	13'h01db: q2 = 16'h0000; // 0x03b6
	13'h01dc: q2 = 16'h8e6c; // 0x03b8
	13'h01dd: q2 = 16'h4a5f; // 0x03ba
	13'h01de: q2 = 16'h33c0; // 0x03bc
	13'h01df: q2 = 16'h0001; // 0x03be
	13'h01e0: q2 = 16'h8070; // 0x03c0
	13'h01e1: q2 = 16'h33ec; // 0x03c2
	13'h01e2: q2 = 16'h0024; // 0x03c4
	13'h01e3: q2 = 16'h0001; // 0x03c6
	13'h01e4: q2 = 16'h8070; // 0x03c8
	13'h01e5: q2 = 16'h6010; // 0x03ca
	13'h01e6: q2 = 16'h3014; // 0x03cc
	13'h01e7: q2 = 16'h48c0; // 0x03ce
	13'h01e8: q2 = 16'h81fc; // 0x03d0
	13'h01e9: q2 = 16'h000a; // 0x03d2
	13'h01ea: q2 = 16'h4840; // 0x03d4
	13'h01eb: q2 = 16'h33c0; // 0x03d6
	13'h01ec: q2 = 16'h0001; // 0x03d8
	13'h01ed: q2 = 16'h8070; // 0x03da
	13'h01ee: q2 = 16'h4246; // 0x03dc
	13'h01ef: q2 = 16'h426e; // 0x03de
	13'h01f0: q2 = 16'hfffa; // 0x03e0
	13'h01f1: q2 = 16'h2a7c; // 0x03e2
	13'h01f2: q2 = 16'h0001; // 0x03e4
	13'h01f3: q2 = 16'h893e; // 0x03e6
	13'h01f4: q2 = 16'h4247; // 0x03e8
	13'h01f5: q2 = 16'hbe79; // 0x03ea
	13'h01f6: q2 = 16'h0001; // 0x03ec
	13'h01f7: q2 = 16'h7fa8; // 0x03ee
	13'h01f8: q2 = 16'h6c00; // 0x03f0
	13'h01f9: q2 = 16'h00fe; // 0x03f2
	13'h01fa: q2 = 16'h3ebc; // 0x03f4
	13'h01fb: q2 = 16'h7700; // 0x03f6
	13'h01fc: q2 = 16'h3f3c; // 0x03f8
	13'h01fd: q2 = 16'h0580; // 0x03fa
	13'h01fe: q2 = 16'h4eb9; // 0x03fc
	13'h01ff: q2 = 16'h0000; // 0x03fe
	13'h0200: q2 = 16'h8e6c; // 0x0400
	13'h0201: q2 = 16'h4a5f; // 0x0402
	13'h0202: q2 = 16'h3d40; // 0x0404
	13'h0203: q2 = 16'hfffe; // 0x0406
	13'h0204: q2 = 16'h3ebc; // 0x0408
	13'h0205: q2 = 16'h6f80; // 0x040a
	13'h0206: q2 = 16'h3f3c; // 0x040c
	13'h0207: q2 = 16'h1800; // 0x040e
	13'h0208: q2 = 16'h4eb9; // 0x0410
	13'h0209: q2 = 16'h0000; // 0x0412
	13'h020a: q2 = 16'h8e6c; // 0x0414
	13'h020b: q2 = 16'h4a5f; // 0x0416
	13'h020c: q2 = 16'h3d40; // 0x0418
	13'h020d: q2 = 16'hfffc; // 0x041a
	13'h020e: q2 = 16'h200e; // 0x041c
	13'h020f: q2 = 16'hd0bc; // 0x041e
	13'h0210: q2 = 16'hffff; // 0x0420
	13'h0211: q2 = 16'hfffc; // 0x0422
	13'h0212: q2 = 16'h2e80; // 0x0424
	13'h0213: q2 = 16'h200e; // 0x0426
	13'h0214: q2 = 16'hd0bc; // 0x0428
	13'h0215: q2 = 16'hffff; // 0x042a
	13'h0216: q2 = 16'hfffe; // 0x042c
	13'h0217: q2 = 16'h2f00; // 0x042e
	13'h0218: q2 = 16'h4eb9; // 0x0430
	13'h0219: q2 = 16'h0000; // 0x0432
	13'h021a: q2 = 16'hbee0; // 0x0434
	13'h021b: q2 = 16'h4a9f; // 0x0436
	13'h021c: q2 = 16'h3ebc; // 0x0438
	13'h021d: q2 = 16'h0001; // 0x043a
	13'h021e: q2 = 16'h3f2e; // 0x043c
	13'h021f: q2 = 16'hfffc; // 0x043e
	13'h0220: q2 = 16'h3f2e; // 0x0440
	13'h0221: q2 = 16'hfffe; // 0x0442
	13'h0222: q2 = 16'h4eb9; // 0x0444
	13'h0223: q2 = 16'h0000; // 0x0446
	13'h0224: q2 = 16'h42d4; // 0x0448
	13'h0225: q2 = 16'h4a9f; // 0x044a
	13'h0226: q2 = 16'h4a40; // 0x044c
	13'h0227: q2 = 16'h66a4; // 0x044e
	13'h0228: q2 = 16'h3ebc; // 0x0450
	13'h0229: q2 = 16'h0001; // 0x0452
	13'h022a: q2 = 16'h3f2e; // 0x0454
	13'h022b: q2 = 16'hfffc; // 0x0456
	13'h022c: q2 = 16'h3f2e; // 0x0458
	13'h022d: q2 = 16'hfffe; // 0x045a
	13'h022e: q2 = 16'h4eb9; // 0x045c
	13'h022f: q2 = 16'h0000; // 0x045e
	13'h0230: q2 = 16'h8744; // 0x0460
	13'h0231: q2 = 16'h4a9f; // 0x0462
	13'h0232: q2 = 16'h4a40; // 0x0464
	13'h0233: q2 = 16'h668c; // 0x0466
	13'h0234: q2 = 16'h3eae; // 0x0468
	13'h0235: q2 = 16'hfffc; // 0x046a
	13'h0236: q2 = 16'h3f2e; // 0x046c
	13'h0237: q2 = 16'hfffe; // 0x046e
	13'h0238: q2 = 16'h4eb9; // 0x0470
	13'h0239: q2 = 16'h0000; // 0x0472
	13'h023a: q2 = 16'h4d7e; // 0x0474
	13'h023b: q2 = 16'h4a5f; // 0x0476
	13'h023c: q2 = 16'h4a40; // 0x0478
	13'h023d: q2 = 16'h6600; // 0x047a
	13'h023e: q2 = 16'hff78; // 0x047c
	13'h023f: q2 = 16'h6004; // 0x047e
	13'h0240: q2 = 16'h6000; // 0x0480
	13'h0241: q2 = 16'hff72; // 0x0482
	13'h0242: q2 = 16'h3aae; // 0x0484
	13'h0243: q2 = 16'hfffe; // 0x0486
	13'h0244: q2 = 16'h3b6e; // 0x0488
	13'h0245: q2 = 16'hfffc; // 0x048a
	13'h0246: q2 = 16'h0002; // 0x048c
	13'h0247: q2 = 16'h3ebc; // 0x048e
	13'h0248: q2 = 16'h0008; // 0x0490
	13'h0249: q2 = 16'h3f3c; // 0x0492
	13'h024a: q2 = 16'h0002; // 0x0494
	13'h024b: q2 = 16'h4eb9; // 0x0496
	13'h024c: q2 = 16'h0000; // 0x0498
	13'h024d: q2 = 16'h8e6c; // 0x049a
	13'h024e: q2 = 16'h4a5f; // 0x049c
	13'h024f: q2 = 16'h3b40; // 0x049e
	13'h0250: q2 = 16'h0006; // 0x04a0
	13'h0251: q2 = 16'hdc6d; // 0x04a2
	13'h0252: q2 = 16'h0006; // 0x04a4
	13'h0253: q2 = 16'h3eb9; // 0x04a6
	13'h0254: q2 = 16'h0001; // 0x04a8
	13'h0255: q2 = 16'h8070; // 0x04aa
	13'h0256: q2 = 16'h4eb9; // 0x04ac
	13'h0257: q2 = 16'h0000; // 0x04ae
	13'h0258: q2 = 16'h3e52; // 0x04b0
	13'h0259: q2 = 16'h3b40; // 0x04b2
	13'h025a: q2 = 16'h0004; // 0x04b4
	13'h025b: q2 = 16'h4a79; // 0x04b6
	13'h025c: q2 = 16'h0001; // 0x04b8
	13'h025d: q2 = 16'h8070; // 0x04ba
	13'h025e: q2 = 16'h6626; // 0x04bc
	13'h025f: q2 = 16'h0c6d; // 0x04be
	13'h0260: q2 = 16'h0005; // 0x04c0
	13'h0261: q2 = 16'h0004; // 0x04c2
	13'h0262: q2 = 16'h6606; // 0x04c4
	13'h0263: q2 = 16'h3d7c; // 0x04c6
	13'h0264: q2 = 16'h0001; // 0x04c8
	13'h0265: q2 = 16'hfffa; // 0x04ca
	13'h0266: q2 = 16'h3039; // 0x04cc
	13'h0267: q2 = 16'h0001; // 0x04ce
	13'h0268: q2 = 16'h7fa8; // 0x04d0
	13'h0269: q2 = 16'h5340; // 0x04d2
	13'h026a: q2 = 16'hb047; // 0x04d4
	13'h026b: q2 = 16'h660c; // 0x04d6
	13'h026c: q2 = 16'h4a6e; // 0x04d8
	13'h026d: q2 = 16'hfffa; // 0x04da
	13'h026e: q2 = 16'h6606; // 0x04dc
	13'h026f: q2 = 16'h3b7c; // 0x04de
	13'h0270: q2 = 16'h0005; // 0x04e0
	13'h0271: q2 = 16'h0004; // 0x04e2
	13'h0272: q2 = 16'hdbfc; // 0x04e4
	13'h0273: q2 = 16'h0000; // 0x04e6
	13'h0274: q2 = 16'h0010; // 0x04e8
	13'h0275: q2 = 16'h5247; // 0x04ea
	13'h0276: q2 = 16'h6000; // 0x04ec
	13'h0277: q2 = 16'hfefc; // 0x04ee
	13'h0278: q2 = 16'h2a7c; // 0x04f0
	13'h0279: q2 = 16'h0001; // 0x04f2
	13'h027a: q2 = 16'h893e; // 0x04f4
	13'h027b: q2 = 16'h4247; // 0x04f6
	13'h027c: q2 = 16'hbc45; // 0x04f8
	13'h027d: q2 = 16'h6740; // 0x04fa
	13'h027e: q2 = 16'hbc45; // 0x04fc
	13'h027f: q2 = 16'h6c10; // 0x04fe
	13'h0280: q2 = 16'h0c6d; // 0x0500
	13'h0281: q2 = 16'h0008; // 0x0502
	13'h0282: q2 = 16'h0006; // 0x0504
	13'h0283: q2 = 16'h6c08; // 0x0506
	13'h0284: q2 = 16'h526d; // 0x0508
	13'h0285: q2 = 16'h0006; // 0x050a
	13'h0286: q2 = 16'h5246; // 0x050c
	13'h0287: q2 = 16'h6012; // 0x050e
	13'h0288: q2 = 16'hbc45; // 0x0510
	13'h0289: q2 = 16'h6f0e; // 0x0512
	13'h028a: q2 = 16'h0c6d; // 0x0514
	13'h028b: q2 = 16'h0002; // 0x0516
	13'h028c: q2 = 16'h0006; // 0x0518
	13'h028d: q2 = 16'h6f06; // 0x051a
	13'h028e: q2 = 16'h536d; // 0x051c
	13'h028f: q2 = 16'h0006; // 0x051e
	13'h0290: q2 = 16'h5346; // 0x0520
	13'h0291: q2 = 16'hdbfc; // 0x0522
	13'h0292: q2 = 16'h0000; // 0x0524
	13'h0293: q2 = 16'h0010; // 0x0526
	13'h0294: q2 = 16'h5247; // 0x0528
	13'h0295: q2 = 16'hbe79; // 0x052a
	13'h0296: q2 = 16'h0001; // 0x052c
	13'h0297: q2 = 16'h7fa8; // 0x052e
	13'h0298: q2 = 16'h6608; // 0x0530
	13'h0299: q2 = 16'h4247; // 0x0532
	13'h029a: q2 = 16'h2a7c; // 0x0534
	13'h029b: q2 = 16'h0001; // 0x0536
	13'h029c: q2 = 16'h893e; // 0x0538
	13'h029d: q2 = 16'h60bc; // 0x053a
	13'h029e: q2 = 16'h2a7c; // 0x053c
	13'h029f: q2 = 16'h0001; // 0x053e
	13'h02a0: q2 = 16'h893e; // 0x0540
	13'h02a1: q2 = 16'h4247; // 0x0542
	13'h02a2: q2 = 16'hbe79; // 0x0544
	13'h02a3: q2 = 16'h0001; // 0x0546
	13'h02a4: q2 = 16'h7fa8; // 0x0548
	13'h02a5: q2 = 16'h6c1a; // 0x054a
	13'h02a6: q2 = 16'h2e8d; // 0x054c
	13'h02a7: q2 = 16'h4eb9; // 0x054e
	13'h02a8: q2 = 16'h0000; // 0x0550
	13'h02a9: q2 = 16'h161a; // 0x0552
	13'h02aa: q2 = 16'h2e8d; // 0x0554
	13'h02ab: q2 = 16'h4eb9; // 0x0556
	13'h02ac: q2 = 16'h0000; // 0x0558
	13'h02ad: q2 = 16'h0f60; // 0x055a
	13'h02ae: q2 = 16'hdbfc; // 0x055c
	13'h02af: q2 = 16'h0000; // 0x055e
	13'h02b0: q2 = 16'h0010; // 0x0560
	13'h02b1: q2 = 16'h5247; // 0x0562
	13'h02b2: q2 = 16'h60de; // 0x0564
	13'h02b3: q2 = 16'h4a9f; // 0x0566
	13'h02b4: q2 = 16'h4cdf; // 0x0568
	13'h02b5: q2 = 16'h30e0; // 0x056a
	13'h02b6: q2 = 16'h4e5e; // 0x056c
	13'h02b7: q2 = 16'h4e75; // 0x056e
	13'h02b8: q2 = 16'h4e56; // 0x0570
	13'h02b9: q2 = 16'hfff2; // 0x0572
	13'h02ba: q2 = 16'h48e7; // 0x0574
	13'h02bb: q2 = 16'h030c; // 0x0576
	13'h02bc: q2 = 16'h4a6e; // 0x0578
	13'h02bd: q2 = 16'h0008; // 0x057a
	13'h02be: q2 = 16'h660a; // 0x057c
	13'h02bf: q2 = 16'h4279; // 0x057e
	13'h02c0: q2 = 16'h0001; // 0x0580
	13'h02c1: q2 = 16'h7fa8; // 0x0582
	13'h02c2: q2 = 16'h6000; // 0x0584
	13'h02c3: q2 = 16'h00f0; // 0x0586
	13'h02c4: q2 = 16'h0c6e; // 0x0588
	13'h02c5: q2 = 16'h0003; // 0x058a
	13'h02c6: q2 = 16'h0008; // 0x058c
	13'h02c7: q2 = 16'h6600; // 0x058e
	13'h02c8: q2 = 16'h00a6; // 0x0590
	13'h02c9: q2 = 16'h33fc; // 0x0592
	13'h02ca: q2 = 16'h0005; // 0x0594
	13'h02cb: q2 = 16'h0001; // 0x0596
	13'h02cc: q2 = 16'h7fa8; // 0x0598
	13'h02cd: q2 = 16'h2a7c; // 0x059a
	13'h02ce: q2 = 16'h0001; // 0x059c
	13'h02cf: q2 = 16'h893e; // 0x059e
	13'h02d0: q2 = 16'h287c; // 0x05a0
	13'h02d1: q2 = 16'h0000; // 0x05a2
	13'h02d2: q2 = 16'hf5cc; // 0x05a4
	13'h02d3: q2 = 16'h4247; // 0x05a6
	13'h02d4: q2 = 16'hbe79; // 0x05a8
	13'h02d5: q2 = 16'h0001; // 0x05aa
	13'h02d6: q2 = 16'h7fa8; // 0x05ac
	13'h02d7: q2 = 16'h6c00; // 0x05ae
	13'h02d8: q2 = 16'h0084; // 0x05b0
	13'h02d9: q2 = 16'h3014; // 0x05b2
	13'h02da: q2 = 16'h4281; // 0x05b4
	13'h02db: q2 = 16'h720a; // 0x05b6
	13'h02dc: q2 = 16'he360; // 0x05b8
	13'h02dd: q2 = 16'h3a80; // 0x05ba
	13'h02de: q2 = 16'h302c; // 0x05bc
	13'h02df: q2 = 16'h0002; // 0x05be
	13'h02e0: q2 = 16'h4281; // 0x05c0
	13'h02e1: q2 = 16'h720a; // 0x05c2
	13'h02e2: q2 = 16'he360; // 0x05c4
	13'h02e3: q2 = 16'h3b40; // 0x05c6
	13'h02e4: q2 = 16'h0002; // 0x05c8
	13'h02e5: q2 = 16'h3b6c; // 0x05ca
	13'h02e6: q2 = 16'h0004; // 0x05cc
	13'h02e7: q2 = 16'h0006; // 0x05ce
	13'h02e8: q2 = 16'h3007; // 0x05d0
	13'h02e9: q2 = 16'h5240; // 0x05d2
	13'h02ea: q2 = 16'h3b40; // 0x05d4
	13'h02eb: q2 = 16'h0004; // 0x05d6
	13'h02ec: q2 = 16'h2e8d; // 0x05d8
	13'h02ed: q2 = 16'h4eb9; // 0x05da
	13'h02ee: q2 = 16'h0000; // 0x05dc
	13'h02ef: q2 = 16'h161a; // 0x05de
	13'h02f0: q2 = 16'h2e8d; // 0x05e0
	13'h02f1: q2 = 16'h4eb9; // 0x05e2
	13'h02f2: q2 = 16'h0000; // 0x05e4
	13'h02f3: q2 = 16'h0f60; // 0x05e6
	13'h02f4: q2 = 16'h3e87; // 0x05e8
	13'h02f5: q2 = 16'h0657; // 0x05ea
	13'h02f6: q2 = 16'h0038; // 0x05ec
	13'h02f7: q2 = 16'h200e; // 0x05ee
	13'h02f8: q2 = 16'hd0bc; // 0x05f0
	13'h02f9: q2 = 16'hffff; // 0x05f2
	13'h02fa: q2 = 16'hfff2; // 0x05f4
	13'h02fb: q2 = 16'h2f00; // 0x05f6
	13'h02fc: q2 = 16'h4eb9; // 0x05f8
	13'h02fd: q2 = 16'h0000; // 0x05fa
	13'h02fe: q2 = 16'h78f6; // 0x05fc
	13'h02ff: q2 = 16'h4a9f; // 0x05fe
	13'h0300: q2 = 16'h3eac; // 0x0600
	13'h0301: q2 = 16'h0006; // 0x0602
	13'h0302: q2 = 16'h4267; // 0x0604
	13'h0303: q2 = 16'h3f2c; // 0x0606
	13'h0304: q2 = 16'h0008; // 0x0608
	13'h0305: q2 = 16'h3f2c; // 0x060a
	13'h0306: q2 = 16'h0002; // 0x060c
	13'h0307: q2 = 16'h200e; // 0x060e
	13'h0308: q2 = 16'hd0bc; // 0x0610
	13'h0309: q2 = 16'hffff; // 0x0612
	13'h030a: q2 = 16'hfff2; // 0x0614
	13'h030b: q2 = 16'h2f00; // 0x0616
	13'h030c: q2 = 16'h4eb9; // 0x0618
	13'h030d: q2 = 16'h0000; // 0x061a
	13'h030e: q2 = 16'h026c; // 0x061c
	13'h030f: q2 = 16'hdefc; // 0x061e
	13'h0310: q2 = 16'h000a; // 0x0620
	13'h0311: q2 = 16'hdbfc; // 0x0622
	13'h0312: q2 = 16'h0000; // 0x0624
	13'h0313: q2 = 16'h0010; // 0x0626
	13'h0314: q2 = 16'hd9fc; // 0x0628
	13'h0315: q2 = 16'h0000; // 0x062a
	13'h0316: q2 = 16'h000a; // 0x062c
	13'h0317: q2 = 16'h5247; // 0x062e
	13'h0318: q2 = 16'h6000; // 0x0630
	13'h0319: q2 = 16'hff76; // 0x0632
	13'h031a: q2 = 16'h6040; // 0x0634
	13'h031b: q2 = 16'h0c6e; // 0x0636
	13'h031c: q2 = 16'h0004; // 0x0638
	13'h031d: q2 = 16'h0008; // 0x063a
	13'h031e: q2 = 16'h6638; // 0x063c
	13'h031f: q2 = 16'h4247; // 0x063e
	13'h0320: q2 = 16'h287c; // 0x0640
	13'h0321: q2 = 16'h0000; // 0x0642
	13'h0322: q2 = 16'hf5cc; // 0x0644
	13'h0323: q2 = 16'hbe79; // 0x0646
	13'h0324: q2 = 16'h0001; // 0x0648
	13'h0325: q2 = 16'h7fa8; // 0x064a
	13'h0326: q2 = 16'h6c28; // 0x064c
	13'h0327: q2 = 16'h4257; // 0x064e
	13'h0328: q2 = 16'h3f3c; // 0x0650
	13'h0329: q2 = 16'h000c; // 0x0652
	13'h032a: q2 = 16'h3f2c; // 0x0654
	13'h032b: q2 = 16'h0008; // 0x0656
	13'h032c: q2 = 16'h3f2c; // 0x0658
	13'h032d: q2 = 16'h0002; // 0x065a
	13'h032e: q2 = 16'h2f3c; // 0x065c
	13'h032f: q2 = 16'h0000; // 0x065e
	13'h0330: q2 = 16'hf5fe; // 0x0660
	13'h0331: q2 = 16'h4eb9; // 0x0662
	13'h0332: q2 = 16'h0000; // 0x0664
	13'h0333: q2 = 16'h026c; // 0x0666
	13'h0334: q2 = 16'hdefc; // 0x0668
	13'h0335: q2 = 16'h000a; // 0x066a
	13'h0336: q2 = 16'h5247; // 0x066c
	13'h0337: q2 = 16'hd9fc; // 0x066e
	13'h0338: q2 = 16'h0000; // 0x0670
	13'h0339: q2 = 16'h000a; // 0x0672
	13'h033a: q2 = 16'h60d0; // 0x0674
	13'h033b: q2 = 16'h4a9f; // 0x0676
	13'h033c: q2 = 16'h4cdf; // 0x0678
	13'h033d: q2 = 16'h3080; // 0x067a
	13'h033e: q2 = 16'h4e5e; // 0x067c
	13'h033f: q2 = 16'h4e75; // 0x067e
	13'h0340: q2 = 16'h4e56; // 0x0680
	13'h0341: q2 = 16'h0000; // 0x0682
	13'h0342: q2 = 16'h48e7; // 0x0684
	13'h0343: q2 = 16'h0104; // 0x0686
	13'h0344: q2 = 16'h33fc; // 0x0688
	13'h0345: q2 = 16'h0001; // 0x068a
	13'h0346: q2 = 16'h0001; // 0x068c
	13'h0347: q2 = 16'h7fa8; // 0x068e
	13'h0348: q2 = 16'h2a7c; // 0x0690
	13'h0349: q2 = 16'h0001; // 0x0692
	13'h034a: q2 = 16'h893e; // 0x0694
	13'h034b: q2 = 16'h3abc; // 0x0696
	13'h034c: q2 = 16'h3c00; // 0x0698
	13'h034d: q2 = 16'h3b7c; // 0x069a
	13'h034e: q2 = 16'h4400; // 0x069c
	13'h034f: q2 = 16'h0002; // 0x069e
	13'h0350: q2 = 16'h3b7c; // 0x06a0
	13'h0351: q2 = 16'h0001; // 0x06a2
	13'h0352: q2 = 16'h0006; // 0x06a4
	13'h0353: q2 = 16'h3b7c; // 0x06a6
	13'h0354: q2 = 16'h0005; // 0x06a8
	13'h0355: q2 = 16'h0004; // 0x06aa
	13'h0356: q2 = 16'h2e8d; // 0x06ac
	13'h0357: q2 = 16'h4eb9; // 0x06ae
	13'h0358: q2 = 16'h0000; // 0x06b0
	13'h0359: q2 = 16'h0f60; // 0x06b2
	13'h035a: q2 = 16'h4a9f; // 0x06b4
	13'h035b: q2 = 16'h4cdf; // 0x06b6
	13'h035c: q2 = 16'h2000; // 0x06b8
	13'h035d: q2 = 16'h4e5e; // 0x06ba
	13'h035e: q2 = 16'h4e75; // 0x06bc
	13'h035f: q2 = 16'h4e56; // 0x06be
	13'h0360: q2 = 16'hfffc; // 0x06c0
	13'h0361: q2 = 16'h48e7; // 0x06c2
	13'h0362: q2 = 16'h0304; // 0x06c4
	13'h0363: q2 = 16'h2a7c; // 0x06c6
	13'h0364: q2 = 16'h0001; // 0x06c8
	13'h0365: q2 = 16'h893e; // 0x06ca
	13'h0366: q2 = 16'h4247; // 0x06cc
	13'h0367: q2 = 16'hbe79; // 0x06ce
	13'h0368: q2 = 16'h0001; // 0x06d0
	13'h0369: q2 = 16'h7fa8; // 0x06d2
	13'h036a: q2 = 16'h6c62; // 0x06d4
	13'h036b: q2 = 16'h4a6d; // 0x06d6
	13'h036c: q2 = 16'h0006; // 0x06d8
	13'h036d: q2 = 16'h6752; // 0x06da
	13'h036e: q2 = 16'h206e; // 0x06dc
	13'h036f: q2 = 16'h0008; // 0x06de
	13'h0370: q2 = 16'h30ad; // 0x06e0
	13'h0371: q2 = 16'h0008; // 0x06e2
	13'h0372: q2 = 16'h206e; // 0x06e4
	13'h0373: q2 = 16'h000c; // 0x06e6
	13'h0374: q2 = 16'h30ad; // 0x06e8
	13'h0375: q2 = 16'h000a; // 0x06ea
	13'h0376: q2 = 16'h2d79; // 0x06ec
	13'h0377: q2 = 16'h0000; // 0x06ee
	13'h0378: q2 = 16'hf600; // 0x06f0
	13'h0379: q2 = 16'hfffc; // 0x06f2
	13'h037a: q2 = 16'h202e; // 0x06f4
	13'h037b: q2 = 16'hfffc; // 0x06f6
	13'h037c: q2 = 16'he780; // 0x06f8
	13'h037d: q2 = 16'h2d40; // 0x06fa
	13'h037e: q2 = 16'hfffc; // 0x06fc
	13'h037f: q2 = 16'h5cae; // 0x06fe
	13'h0380: q2 = 16'hfffc; // 0x0700
	13'h0381: q2 = 16'h206e; // 0x0702
	13'h0382: q2 = 16'hfffc; // 0x0704
	13'h0383: q2 = 16'h3010; // 0x0706
	13'h0384: q2 = 16'hc07c; // 0x0708
	13'h0385: q2 = 16'h0ff0; // 0x070a
	13'h0386: q2 = 16'hb07c; // 0x070c
	13'h0387: q2 = 16'h0950; // 0x070e
	13'h0388: q2 = 16'h6610; // 0x0710
	13'h0389: q2 = 16'h206e; // 0x0712
	13'h038a: q2 = 16'hfffc; // 0x0714
	13'h038b: q2 = 16'h3010; // 0x0716
	13'h038c: q2 = 16'hc07c; // 0x0718
	13'h038d: q2 = 16'hf00f; // 0x071a
	13'h038e: q2 = 16'hb07c; // 0x071c
	13'h038f: q2 = 16'h2002; // 0x071e
	13'h0390: q2 = 16'h6708; // 0x0720
	13'h0391: q2 = 16'h33fc; // 0x0722
	13'h0392: q2 = 16'h0001; // 0x0724
	13'h0393: q2 = 16'h0001; // 0x0726
	13'h0394: q2 = 16'h75e6; // 0x0728
	13'h0395: q2 = 16'h7001; // 0x072a
	13'h0396: q2 = 16'h600c; // 0x072c
	13'h0397: q2 = 16'hdbfc; // 0x072e
	13'h0398: q2 = 16'h0000; // 0x0730
	13'h0399: q2 = 16'h0010; // 0x0732
	13'h039a: q2 = 16'h5247; // 0x0734
	13'h039b: q2 = 16'h6096; // 0x0736
	13'h039c: q2 = 16'h4240; // 0x0738
	13'h039d: q2 = 16'h4a9f; // 0x073a
	13'h039e: q2 = 16'h4cdf; // 0x073c
	13'h039f: q2 = 16'h2080; // 0x073e
	13'h03a0: q2 = 16'h4e5e; // 0x0740
	13'h03a1: q2 = 16'h4e75; // 0x0742
	13'h03a2: q2 = 16'h4e56; // 0x0744
	13'h03a3: q2 = 16'h0000; // 0x0746
	13'h03a4: q2 = 16'h48e7; // 0x0748
	13'h03a5: q2 = 16'h3f04; // 0x074a
	13'h03a6: q2 = 16'h2a7c; // 0x074c
	13'h03a7: q2 = 16'h0001; // 0x074e
	13'h03a8: q2 = 16'h893e; // 0x0750
	13'h03a9: q2 = 16'h4247; // 0x0752
	13'h03aa: q2 = 16'hbe79; // 0x0754
	13'h03ab: q2 = 16'h0001; // 0x0756
	13'h03ac: q2 = 16'h7fa8; // 0x0758
	13'h03ad: q2 = 16'h6c60; // 0x075a
	13'h03ae: q2 = 16'h4a6d; // 0x075c
	13'h03af: q2 = 16'h0006; // 0x075e
	13'h03b0: q2 = 16'h6750; // 0x0760
	13'h03b1: q2 = 16'h4a6e; // 0x0762
	13'h03b2: q2 = 16'h000c; // 0x0764
	13'h03b3: q2 = 16'h6710; // 0x0766
	13'h03b4: q2 = 16'h3c15; // 0x0768
	13'h03b5: q2 = 16'h3a2d; // 0x076a
	13'h03b6: q2 = 16'h0002; // 0x076c
	13'h03b7: q2 = 16'h383c; // 0x076e
	13'h03b8: q2 = 16'h1000; // 0x0770
	13'h03b9: q2 = 16'h363c; // 0x0772
	13'h03ba: q2 = 16'h1000; // 0x0774
	13'h03bb: q2 = 16'h6010; // 0x0776
	13'h03bc: q2 = 16'h3c2d; // 0x0778
	13'h03bd: q2 = 16'h0008; // 0x077a
	13'h03be: q2 = 16'h3a2d; // 0x077c
	13'h03bf: q2 = 16'h000a; // 0x077e
	13'h03c0: q2 = 16'h382d; // 0x0780
	13'h03c1: q2 = 16'h000c; // 0x0782
	13'h03c2: q2 = 16'h362d; // 0x0784
	13'h03c3: q2 = 16'h000e; // 0x0786
	13'h03c4: q2 = 16'h3eae; // 0x0788
	13'h03c5: q2 = 16'h0008; // 0x078a
	13'h03c6: q2 = 16'h3006; // 0x078c
	13'h03c7: q2 = 16'h9157; // 0x078e
	13'h03c8: q2 = 16'h4eb9; // 0x0790
	13'h03c9: q2 = 16'h0000; // 0x0792
	13'h03ca: q2 = 16'h09a2; // 0x0794
	13'h03cb: q2 = 16'hb044; // 0x0796
	13'h03cc: q2 = 16'h6c18; // 0x0798
	13'h03cd: q2 = 16'h3eae; // 0x079a
	13'h03ce: q2 = 16'h000a; // 0x079c
	13'h03cf: q2 = 16'h3005; // 0x079e
	13'h03d0: q2 = 16'h9157; // 0x07a0
	13'h03d1: q2 = 16'h4eb9; // 0x07a2
	13'h03d2: q2 = 16'h0000; // 0x07a4
	13'h03d3: q2 = 16'h09a2; // 0x07a6
	13'h03d4: q2 = 16'hb043; // 0x07a8
	13'h03d5: q2 = 16'h6c06; // 0x07aa
	13'h03d6: q2 = 16'h3007; // 0x07ac
	13'h03d7: q2 = 16'h5240; // 0x07ae
	13'h03d8: q2 = 16'h600c; // 0x07b0
	13'h03d9: q2 = 16'hdbfc; // 0x07b2
	13'h03da: q2 = 16'h0000; // 0x07b4
	13'h03db: q2 = 16'h0010; // 0x07b6
	13'h03dc: q2 = 16'h5247; // 0x07b8
	13'h03dd: q2 = 16'h6098; // 0x07ba
	13'h03de: q2 = 16'h4240; // 0x07bc
	13'h03df: q2 = 16'h4a9f; // 0x07be
	13'h03e0: q2 = 16'h4cdf; // 0x07c0
	13'h03e1: q2 = 16'h20f8; // 0x07c2
	13'h03e2: q2 = 16'h4e5e; // 0x07c4
	13'h03e3: q2 = 16'h4e75; // 0x07c6
	13'h03e4: q2 = 16'h4e56; // 0x07c8
	13'h03e5: q2 = 16'h0000; // 0x07ca
	13'h03e6: q2 = 16'h48e7; // 0x07cc
	13'h03e7: q2 = 16'h0304; // 0x07ce
	13'h03e8: q2 = 16'h4247; // 0x07d0
	13'h03e9: q2 = 16'h2a7c; // 0x07d2
	13'h03ea: q2 = 16'h0001; // 0x07d4
	13'h03eb: q2 = 16'h8628; // 0x07d6
	13'h03ec: q2 = 16'hbe7c; // 0x07d8
	13'h03ed: q2 = 16'h0001; // 0x07da
	13'h03ee: q2 = 16'h6e46; // 0x07dc
	13'h03ef: q2 = 16'h42ad; // 0x07de
	13'h03f0: q2 = 16'h0004; // 0x07e0
	13'h03f1: q2 = 16'h4a79; // 0x07e2
	13'h03f2: q2 = 16'h0001; // 0x07e4
	13'h03f3: q2 = 16'h7580; // 0x07e6
	13'h03f4: q2 = 16'h6f0c; // 0x07e8
	13'h03f5: q2 = 16'h3079; // 0x07ea
	13'h03f6: q2 = 16'h0001; // 0x07ec
	13'h03f7: q2 = 16'h7580; // 0x07ee
	13'h03f8: q2 = 16'h2b48; // 0x07f0
	13'h03f9: q2 = 16'h0018; // 0x07f2
	13'h03fa: q2 = 16'h600a; // 0x07f4
	13'h03fb: q2 = 16'h3079; // 0x07f6
	13'h03fc: q2 = 16'h0001; // 0x07f8
	13'h03fd: q2 = 16'h7582; // 0x07fa
	13'h03fe: q2 = 16'h2b48; // 0x07fc
	13'h03ff: q2 = 16'h0018; // 0x07fe
	13'h0400: q2 = 16'h3b79; // 0x0800
	13'h0401: q2 = 16'h0001; // 0x0802
	13'h0402: q2 = 16'h757a; // 0x0804
	13'h0403: q2 = 16'h0002; // 0x0806
	13'h0404: q2 = 16'h426d; // 0x0808
	13'h0405: q2 = 16'h001e; // 0x080a
	13'h0406: q2 = 16'h426d; // 0x080c
	13'h0407: q2 = 16'h0020; // 0x080e
	13'h0408: q2 = 16'h3b7c; // 0x0810
	13'h0409: q2 = 16'h0001; // 0x0812
	13'h040a: q2 = 16'h0022; // 0x0814
	13'h040b: q2 = 16'h426d; // 0x0816
	13'h040c: q2 = 16'h0024; // 0x0818
	13'h040d: q2 = 16'h5247; // 0x081a
	13'h040e: q2 = 16'hdbfc; // 0x081c
	13'h040f: q2 = 16'h0000; // 0x081e
	13'h0410: q2 = 16'h0026; // 0x0820
	13'h0411: q2 = 16'h60b4; // 0x0822
	13'h0412: q2 = 16'h2ebc; // 0x0824
	13'h0413: q2 = 16'h0000; // 0x0826
	13'h0414: q2 = 16'hf76e; // 0x0828
	13'h0415: q2 = 16'h2f3c; // 0x082a
	13'h0416: q2 = 16'h0001; // 0x082c
	13'h0417: q2 = 16'h8630; // 0x082e
	13'h0418: q2 = 16'h4eb9; // 0x0830
	13'h0419: q2 = 16'h0000; // 0x0832
	13'h041a: q2 = 16'h0750; // 0x0834
	13'h041b: q2 = 16'h4a9f; // 0x0836
	13'h041c: q2 = 16'h2ebc; // 0x0838
	13'h041d: q2 = 16'h0000; // 0x083a
	13'h041e: q2 = 16'hf772; // 0x083c
	13'h041f: q2 = 16'h2f3c; // 0x083e
	13'h0420: q2 = 16'h0001; // 0x0840
	13'h0421: q2 = 16'h8656; // 0x0842
	13'h0422: q2 = 16'h4eb9; // 0x0844
	13'h0423: q2 = 16'h0000; // 0x0846
	13'h0424: q2 = 16'h0750; // 0x0848
	13'h0425: q2 = 16'h4a9f; // 0x084a
	13'h0426: q2 = 16'h4a9f; // 0x084c
	13'h0427: q2 = 16'h4cdf; // 0x084e
	13'h0428: q2 = 16'h2080; // 0x0850
	13'h0429: q2 = 16'h4e5e; // 0x0852
	13'h042a: q2 = 16'h4e75; // 0x0854
	13'h042b: q2 = 16'h4e56; // 0x0856
	13'h042c: q2 = 16'hffee; // 0x0858
	13'h042d: q2 = 16'h3ebc; // 0x085a
	13'h042e: q2 = 16'h001a; // 0x085c
	13'h042f: q2 = 16'h4eb9; // 0x085e
	13'h0430: q2 = 16'h0000; // 0x0860
	13'h0431: q2 = 16'h8a22; // 0x0862
	13'h0432: q2 = 16'h3ebc; // 0x0864
	13'h0433: q2 = 16'h0037; // 0x0866
	13'h0434: q2 = 16'h200e; // 0x0868
	13'h0435: q2 = 16'hd0bc; // 0x086a
	13'h0436: q2 = 16'hffff; // 0x086c
	13'h0437: q2 = 16'hfff2; // 0x086e
	13'h0438: q2 = 16'h2f00; // 0x0870
	13'h0439: q2 = 16'h4eb9; // 0x0872
	13'h043a: q2 = 16'h0000; // 0x0874
	13'h043b: q2 = 16'h78f6; // 0x0876
	13'h043c: q2 = 16'h4a9f; // 0x0878
	13'h043d: q2 = 16'h200e; // 0x087a
	13'h043e: q2 = 16'hd0bc; // 0x087c
	13'h043f: q2 = 16'hffff; // 0x087e
	13'h0440: q2 = 16'hfff2; // 0x0880
	13'h0441: q2 = 16'h2e80; // 0x0882
	13'h0442: q2 = 16'h3f2e; // 0x0884
	13'h0443: q2 = 16'h0008; // 0x0886
	13'h0444: q2 = 16'h4eb9; // 0x0888
	13'h0445: q2 = 16'h0000; // 0x088a
	13'h0446: q2 = 16'h0798; // 0x088c
	13'h0447: q2 = 16'h4a5f; // 0x088e
	13'h0448: q2 = 16'h3ebc; // 0x0890
	13'h0449: q2 = 16'h003e; // 0x0892
	13'h044a: q2 = 16'h4267; // 0x0894
	13'h044b: q2 = 16'h3f3c; // 0x0896
	13'h044c: q2 = 16'h0064; // 0x0898
	13'h044d: q2 = 16'h3f3c; // 0x089a
	13'h044e: q2 = 16'h0010; // 0x089c
	13'h044f: q2 = 16'h200e; // 0x089e
	13'h0450: q2 = 16'hd0bc; // 0x08a0
	13'h0451: q2 = 16'hffff; // 0x08a2
	13'h0452: q2 = 16'hfff2; // 0x08a4
	13'h0453: q2 = 16'h2f00; // 0x08a6
	13'h0454: q2 = 16'h4eb9; // 0x08a8
	13'h0455: q2 = 16'h0000; // 0x08aa
	13'h0456: q2 = 16'h026c; // 0x08ac
	13'h0457: q2 = 16'hdefc; // 0x08ae
	13'h0458: q2 = 16'h000a; // 0x08b0
	13'h0459: q2 = 16'h2eb9; // 0x08b2
	13'h045a: q2 = 16'h0000; // 0x08b4
	13'h045b: q2 = 16'hf774; // 0x08b6
	13'h045c: q2 = 16'h4eb9; // 0x08b8
	13'h045d: q2 = 16'h0000; // 0x08ba
	13'h045e: q2 = 16'h3da4; // 0x08bc
	13'h045f: q2 = 16'h3ebc; // 0x08be
	13'h0460: q2 = 16'h0001; // 0x08c0
	13'h0461: q2 = 16'h3f3c; // 0x08c2
	13'h0462: q2 = 16'h0018; // 0x08c4
	13'h0463: q2 = 16'h3f3c; // 0x08c6
	13'h0464: q2 = 16'h0064; // 0x08c8
	13'h0465: q2 = 16'h3f3c; // 0x08ca
	13'h0466: q2 = 16'h0012; // 0x08cc
	13'h0467: q2 = 16'h2f3c; // 0x08ce
	13'h0468: q2 = 16'h0000; // 0x08d0
	13'h0469: q2 = 16'hf778; // 0x08d2
	13'h046a: q2 = 16'h4eb9; // 0x08d4
	13'h046b: q2 = 16'h0000; // 0x08d6
	13'h046c: q2 = 16'h026c; // 0x08d8
	13'h046d: q2 = 16'hdefc; // 0x08da
	13'h046e: q2 = 16'h000a; // 0x08dc
	13'h046f: q2 = 16'h3ebc; // 0x08de
	13'h0470: q2 = 16'h0001; // 0x08e0
	13'h0471: q2 = 16'h3f3c; // 0x08e2
	13'h0472: q2 = 16'h0009; // 0x08e4
	13'h0473: q2 = 16'h3f3c; // 0x08e6
	13'h0474: q2 = 16'h0064; // 0x08e8
	13'h0475: q2 = 16'h3f3c; // 0x08ea
	13'h0476: q2 = 16'h0010; // 0x08ec
	13'h0477: q2 = 16'h2f3c; // 0x08ee
	13'h0478: q2 = 16'h0000; // 0x08f0
	13'h0479: q2 = 16'hf779; // 0x08f2
	13'h047a: q2 = 16'h4eb9; // 0x08f4
	13'h047b: q2 = 16'h0000; // 0x08f6
	13'h047c: q2 = 16'h026c; // 0x08f8
	13'h047d: q2 = 16'hdefc; // 0x08fa
	13'h047e: q2 = 16'h000a; // 0x08fc
	13'h047f: q2 = 16'h4e5e; // 0x08fe
	13'h0480: q2 = 16'h4e75; // 0x0900
	13'h0481: q2 = 16'h4e56; // 0x0902
	13'h0482: q2 = 16'hfffc; // 0x0904
	13'h0483: q2 = 16'h2eb9; // 0x0906
	13'h0484: q2 = 16'h0000; // 0x0908
	13'h0485: q2 = 16'hf51c; // 0x090a
	13'h0486: q2 = 16'h6132; // 0x090c
	13'h0487: q2 = 16'h2039; // 0x090e
	13'h0488: q2 = 16'h0000; // 0x0910
	13'h0489: q2 = 16'hf51c; // 0x0912
	13'h048a: q2 = 16'hd0b9; // 0x0914
	13'h048b: q2 = 16'h0000; // 0x0916
	13'h048c: q2 = 16'hf520; // 0x0918
	13'h048d: q2 = 16'h2e80; // 0x091a
	13'h048e: q2 = 16'h6122; // 0x091c
	13'h048f: q2 = 16'h2039; // 0x091e
	13'h0490: q2 = 16'h0000; // 0x0920
	13'h0491: q2 = 16'hf520; // 0x0922
	13'h0492: q2 = 16'he380; // 0x0924
	13'h0493: q2 = 16'hd0b9; // 0x0926
	13'h0494: q2 = 16'h0000; // 0x0928
	13'h0495: q2 = 16'hf51c; // 0x092a
	13'h0496: q2 = 16'h2e80; // 0x092c
	13'h0497: q2 = 16'h6110; // 0x092e
	13'h0498: q2 = 16'h4eb9; // 0x0930
	13'h0499: q2 = 16'h0000; // 0x0932
	13'h049a: q2 = 16'hb366; // 0x0934
	13'h049b: q2 = 16'h4eb9; // 0x0936
	13'h049c: q2 = 16'h0000; // 0x0938
	13'h049d: q2 = 16'hba28; // 0x093a
	13'h049e: q2 = 16'h4e5e; // 0x093c
	13'h049f: q2 = 16'h4e75; // 0x093e
	13'h04a0: q2 = 16'h4e56; // 0x0940
	13'h04a1: q2 = 16'hfff8; // 0x0942
	13'h04a2: q2 = 16'h426e; // 0x0944
	13'h04a3: q2 = 16'hfffc; // 0x0946
	13'h04a4: q2 = 16'h426e; // 0x0948
	13'h04a5: q2 = 16'hfffe; // 0x094a
	13'h04a6: q2 = 16'h0c6e; // 0x094c
	13'h04a7: q2 = 16'h0010; // 0x094e
	13'h04a8: q2 = 16'hfffe; // 0x0950
	13'h04a9: q2 = 16'h6c18; // 0x0952
	13'h04aa: q2 = 16'h302e; // 0x0954
	13'h04ab: q2 = 16'hfffe; // 0x0956
	13'h04ac: q2 = 16'he340; // 0x0958
	13'h04ad: q2 = 16'h48c0; // 0x095a
	13'h04ae: q2 = 16'hd0ae; // 0x095c
	13'h04af: q2 = 16'h0008; // 0x095e
	13'h04b0: q2 = 16'h2040; // 0x0960
	13'h04b1: q2 = 16'h30ae; // 0x0962
	13'h04b2: q2 = 16'hfffc; // 0x0964
	13'h04b3: q2 = 16'h526e; // 0x0966
	13'h04b4: q2 = 16'hfffe; // 0x0968
	13'h04b5: q2 = 16'h60e0; // 0x096a
	13'h04b6: q2 = 16'h206e; // 0x096c
	13'h04b7: q2 = 16'h0008; // 0x096e
	13'h04b8: q2 = 16'h317c; // 0x0970
	13'h04b9: q2 = 16'h0083; // 0x0972
	13'h04ba: q2 = 16'h001e; // 0x0974
	13'h04bb: q2 = 16'h4e5e; // 0x0976
	13'h04bc: q2 = 16'h4e75; // 0x0978
	13'h04bd: q2 = 16'h4e56; // 0x097a
	13'h04be: q2 = 16'hfffc; // 0x097c
	13'h04bf: q2 = 16'h48e7; // 0x097e
	13'h04c0: q2 = 16'h0304; // 0x0980
	13'h04c1: q2 = 16'h4eb9; // 0x0982
	13'h04c2: q2 = 16'h0000; // 0x0984
	13'h04c3: q2 = 16'h8902; // 0x0986
	13'h04c4: q2 = 16'h4eb9; // 0x0988
	13'h04c5: q2 = 16'h0000; // 0x098a
	13'h04c6: q2 = 16'h8ea8; // 0x098c
	13'h04c7: q2 = 16'h4eb9; // 0x098e
	13'h04c8: q2 = 16'h0000; // 0x0990
	13'h04c9: q2 = 16'h0fd4; // 0x0992
	13'h04ca: q2 = 16'h23fc; // 0x0994
	13'h04cb: q2 = 16'h0000; // 0x0996
	13'h04cc: q2 = 16'h0001; // 0x0998
	13'h04cd: q2 = 16'h0001; // 0x099a
	13'h04ce: q2 = 16'h7596; // 0x099c
	13'h04cf: q2 = 16'h4247; // 0x099e
	13'h04d0: q2 = 16'h2a7c; // 0x09a0
	13'h04d1: q2 = 16'h0001; // 0x09a2
	13'h04d2: q2 = 16'h86dc; // 0x09a4
	13'h04d3: q2 = 16'hbe7c; // 0x09a6
	13'h04d4: q2 = 16'h0030; // 0x09a8
	13'h04d5: q2 = 16'h6c14; // 0x09aa
	13'h04d6: q2 = 16'h4215; // 0x09ac
	13'h04d7: q2 = 16'h422d; // 0x09ae
	13'h04d8: q2 = 16'h0001; // 0x09b0
	13'h04d9: q2 = 16'h422d; // 0x09b2
	13'h04da: q2 = 16'h0002; // 0x09b4
	13'h04db: q2 = 16'h422d; // 0x09b6
	13'h04dc: q2 = 16'h0003; // 0x09b8
	13'h04dd: q2 = 16'h5247; // 0x09ba
	13'h04de: q2 = 16'h588d; // 0x09bc
	13'h04df: q2 = 16'h60e6; // 0x09be
	13'h04e0: q2 = 16'h4240; // 0x09c0
	13'h04e1: q2 = 16'h33c0; // 0x09c2
	13'h04e2: q2 = 16'h0001; // 0x09c4
	13'h04e3: q2 = 16'h86aa; // 0x09c6
	13'h04e4: q2 = 16'h33c0; // 0x09c8
	13'h04e5: q2 = 16'h0001; // 0x09ca
	13'h04e6: q2 = 16'h8680; // 0x09cc
	13'h04e7: q2 = 16'h4279; // 0x09ce
	13'h04e8: q2 = 16'h0001; // 0x09d0
	13'h04e9: q2 = 16'h7fcc; // 0x09d2
	13'h04ea: q2 = 16'h4279; // 0x09d4
	13'h04eb: q2 = 16'h0001; // 0x09d6
	13'h04ec: q2 = 16'h7fa6; // 0x09d8
	13'h04ed: q2 = 16'h4279; // 0x09da
	13'h04ee: q2 = 16'h0001; // 0x09dc
	13'h04ef: q2 = 16'h8052; // 0x09de
	13'h04f0: q2 = 16'h33fc; // 0x09e0
	13'h04f1: q2 = 16'h0001; // 0x09e2
	13'h04f2: q2 = 16'h0001; // 0x09e4
	13'h04f3: q2 = 16'h757c; // 0x09e6
	13'h04f4: q2 = 16'h4279; // 0x09e8
	13'h04f5: q2 = 16'h0001; // 0x09ea
	13'h04f6: q2 = 16'h7fa8; // 0x09ec
	13'h04f7: q2 = 16'h33fc; // 0x09ee
	13'h04f8: q2 = 16'h0001; // 0x09f0
	13'h04f9: q2 = 16'h0001; // 0x09f2
	13'h04fa: q2 = 16'h805a; // 0x09f4
	13'h04fb: q2 = 16'h4eb9; // 0x09f6
	13'h04fc: q2 = 16'h0000; // 0x09f8
	13'h04fd: q2 = 16'h209c; // 0x09fa
	13'h04fe: q2 = 16'h2d79; // 0x09fc
	13'h04ff: q2 = 16'h0000; // 0x09fe
	13'h0500: q2 = 16'hf77a; // 0x0a00
	13'h0501: q2 = 16'hfffc; // 0x0a02
	13'h0502: q2 = 16'h206e; // 0x0a04
	13'h0503: q2 = 16'hfffc; // 0x0a06
	13'h0504: q2 = 16'h317c; // 0x0a08
	13'h0505: q2 = 16'h0003; // 0x0a0a
	13'h0506: q2 = 16'h001e; // 0x0a0c
	13'h0507: q2 = 16'h206e; // 0x0a0e
	13'h0508: q2 = 16'hfffc; // 0x0a10
	13'h0509: q2 = 16'h317c; // 0x0a12
	13'h050a: q2 = 16'h0007; // 0x0a14
	13'h050b: q2 = 16'h0016; // 0x0a16
	13'h050c: q2 = 16'h4a9f; // 0x0a18
	13'h050d: q2 = 16'h4cdf; // 0x0a1a
	13'h050e: q2 = 16'h2080; // 0x0a1c
	13'h050f: q2 = 16'h4e5e; // 0x0a1e
	13'h0510: q2 = 16'h4e75; // 0x0a20
	13'h0511: q2 = 16'h4e56; // 0x0a22
	13'h0512: q2 = 16'hffde; // 0x0a24
	13'h0513: q2 = 16'h48e7; // 0x0a26
	13'h0514: q2 = 16'h0104; // 0x0a28
	13'h0515: q2 = 16'h302e; // 0x0a2a
	13'h0516: q2 = 16'h0008; // 0x0a2c
	13'h0517: q2 = 16'hc1fc; // 0x0a2e
	13'h0518: q2 = 16'h0005; // 0x0a30
	13'h0519: q2 = 16'h48c0; // 0x0a32
	13'h051a: q2 = 16'h2a40; // 0x0a34
	13'h051b: q2 = 16'hdbfc; // 0x0a36
	13'h051c: q2 = 16'h0000; // 0x0a38
	13'h051d: q2 = 16'hf77e; // 0x0a3a
	13'h051e: q2 = 16'h1015; // 0x0a3c
	13'h051f: q2 = 16'h4880; // 0x0a3e
	13'h0520: q2 = 16'h3e80; // 0x0a40
	13'h0521: q2 = 16'h200e; // 0x0a42
	13'h0522: q2 = 16'hd0bc; // 0x0a44
	13'h0523: q2 = 16'hffff; // 0x0a46
	13'h0524: q2 = 16'hffde; // 0x0a48
	13'h0525: q2 = 16'h2f00; // 0x0a4a
	13'h0526: q2 = 16'h4eb9; // 0x0a4c
	13'h0527: q2 = 16'h0000; // 0x0a4e
	13'h0528: q2 = 16'h78f6; // 0x0a50
	13'h0529: q2 = 16'h4a9f; // 0x0a52
	13'h052a: q2 = 16'h102d; // 0x0a54
	13'h052b: q2 = 16'h0004; // 0x0a56
	13'h052c: q2 = 16'h4880; // 0x0a58
	13'h052d: q2 = 16'h3e80; // 0x0a5a
	13'h052e: q2 = 16'h102d; // 0x0a5c
	13'h052f: q2 = 16'h0003; // 0x0a5e
	13'h0530: q2 = 16'h4880; // 0x0a60
	13'h0531: q2 = 16'h3f00; // 0x0a62
	13'h0532: q2 = 16'h102d; // 0x0a64
	13'h0533: q2 = 16'h0002; // 0x0a66
	13'h0534: q2 = 16'h4880; // 0x0a68
	13'h0535: q2 = 16'h3f00; // 0x0a6a
	13'h0536: q2 = 16'h102d; // 0x0a6c
	13'h0537: q2 = 16'h0001; // 0x0a6e
	13'h0538: q2 = 16'h4880; // 0x0a70
	13'h0539: q2 = 16'h3f00; // 0x0a72
	13'h053a: q2 = 16'h200e; // 0x0a74
	13'h053b: q2 = 16'hd0bc; // 0x0a76
	13'h053c: q2 = 16'hffff; // 0x0a78
	13'h053d: q2 = 16'hffde; // 0x0a7a
	13'h053e: q2 = 16'h2f00; // 0x0a7c
	13'h053f: q2 = 16'h4eb9; // 0x0a7e
	13'h0540: q2 = 16'h0000; // 0x0a80
	13'h0541: q2 = 16'h026c; // 0x0a82
	13'h0542: q2 = 16'hdefc; // 0x0a84
	13'h0543: q2 = 16'h000a; // 0x0a86
	13'h0544: q2 = 16'h4a9f; // 0x0a88
	13'h0545: q2 = 16'h4cdf; // 0x0a8a
	13'h0546: q2 = 16'h2000; // 0x0a8c
	13'h0547: q2 = 16'h4e5e; // 0x0a8e
	13'h0548: q2 = 16'h4e75; // 0x0a90
	13'h0549: q2 = 16'h4e56; // 0x0a92
	13'h054a: q2 = 16'hffee; // 0x0a94
	13'h054b: q2 = 16'h48e7; // 0x0a96
	13'h054c: q2 = 16'h1f1c; // 0x0a98
	13'h054d: q2 = 16'h287c; // 0x0a9a
	13'h054e: q2 = 16'h0001; // 0x0a9c
	13'h054f: q2 = 16'h8628; // 0x0a9e
	13'h0550: q2 = 16'h267c; // 0x0aa0
	13'h0551: q2 = 16'h0001; // 0x0aa2
	13'h0552: q2 = 16'h864e; // 0x0aa4
	13'h0553: q2 = 16'h4a79; // 0x0aa6
	13'h0554: q2 = 16'h0001; // 0x0aa8
	13'h0555: q2 = 16'h7fc6; // 0x0aaa
	13'h0556: q2 = 16'h6608; // 0x0aac
	13'h0557: q2 = 16'h4a79; // 0x0aae
	13'h0558: q2 = 16'h0001; // 0x0ab0
	13'h0559: q2 = 16'h8054; // 0x0ab2
	13'h055a: q2 = 16'h6608; // 0x0ab4
	13'h055b: q2 = 16'h3d7c; // 0x0ab6
	13'h055c: q2 = 16'h0025; // 0x0ab8
	13'h055d: q2 = 16'hffee; // 0x0aba
	13'h055e: q2 = 16'h6006; // 0x0abc
	13'h055f: q2 = 16'h3d7c; // 0x0abe
	13'h0560: q2 = 16'h0027; // 0x0ac0
	13'h0561: q2 = 16'hffee; // 0x0ac2
	13'h0562: q2 = 16'h3eae; // 0x0ac4
	13'h0563: q2 = 16'hffee; // 0x0ac6
	13'h0564: q2 = 16'h4267; // 0x0ac8
	13'h0565: q2 = 16'h4267; // 0x0aca
	13'h0566: q2 = 16'h3f3c; // 0x0acc
	13'h0567: q2 = 16'h001f; // 0x0ace
	13'h0568: q2 = 16'h200c; // 0x0ad0
	13'h0569: q2 = 16'h5080; // 0x0ad2
	13'h056a: q2 = 16'h2f00; // 0x0ad4
	13'h056b: q2 = 16'h4eb9; // 0x0ad6
	13'h056c: q2 = 16'h0000; // 0x0ad8
	13'h056d: q2 = 16'h026c; // 0x0ada
	13'h056e: q2 = 16'hdefc; // 0x0adc
	13'h056f: q2 = 16'h000a; // 0x0ade
	13'h0570: q2 = 16'h200c; // 0x0ae0
	13'h0571: q2 = 16'h5080; // 0x0ae2
	13'h0572: q2 = 16'h2e80; // 0x0ae4
	13'h0573: q2 = 16'h4eb9; // 0x0ae6
	13'h0574: q2 = 16'h0000; // 0x0ae8
	13'h0575: q2 = 16'h072e; // 0x0aea
	13'h0576: q2 = 16'h3c00; // 0x0aec
	13'h0577: q2 = 16'h3006; // 0x0aee
	13'h0578: q2 = 16'h5740; // 0x0af0
	13'h0579: q2 = 16'h4281; // 0x0af2
	13'h057a: q2 = 16'h720a; // 0x0af4
	13'h057b: q2 = 16'he360; // 0x0af6
	13'h057c: q2 = 16'h3940; // 0x0af8
	13'h057d: q2 = 16'h0014; // 0x0afa
	13'h057e: q2 = 16'h4245; // 0x0afc
	13'h057f: q2 = 16'h0c79; // 0x0afe
	13'h0580: q2 = 16'h0002; // 0x0b00
	13'h0581: q2 = 16'h0001; // 0x0b02
	13'h0582: q2 = 16'h87dc; // 0x0b04
	13'h0583: q2 = 16'h664c; // 0x0b06
	13'h0584: q2 = 16'h4a79; // 0x0b08
	13'h0585: q2 = 16'h0001; // 0x0b0a
	13'h0586: q2 = 16'h7fc6; // 0x0b0c
	13'h0587: q2 = 16'h660a; // 0x0b0e
	13'h0588: q2 = 16'h0c79; // 0x0b10
	13'h0589: q2 = 16'h0001; // 0x0b12
	13'h058a: q2 = 16'h0001; // 0x0b14
	13'h058b: q2 = 16'h8054; // 0x0b16
	13'h058c: q2 = 16'h6608; // 0x0b18
	13'h058d: q2 = 16'h3d7c; // 0x0b1a
	13'h058e: q2 = 16'h0025; // 0x0b1c
	13'h058f: q2 = 16'hffee; // 0x0b1e
	13'h0590: q2 = 16'h6006; // 0x0b20
	13'h0591: q2 = 16'h3d7c; // 0x0b22
	13'h0592: q2 = 16'h0027; // 0x0b24
	13'h0593: q2 = 16'hffee; // 0x0b26
	13'h0594: q2 = 16'h3eae; // 0x0b28
	13'h0595: q2 = 16'hffee; // 0x0b2a
	13'h0596: q2 = 16'h4267; // 0x0b2c
	13'h0597: q2 = 16'h3f3c; // 0x0b2e
	13'h0598: q2 = 16'hffe1; // 0x0b30
	13'h0599: q2 = 16'h3f3c; // 0x0b32
	13'h059a: q2 = 16'h001f; // 0x0b34
	13'h059b: q2 = 16'h200b; // 0x0b36
	13'h059c: q2 = 16'h5080; // 0x0b38
	13'h059d: q2 = 16'h2f00; // 0x0b3a
	13'h059e: q2 = 16'h4eb9; // 0x0b3c
	13'h059f: q2 = 16'h0000; // 0x0b3e
	13'h05a0: q2 = 16'h026c; // 0x0b40
	13'h05a1: q2 = 16'hdefc; // 0x0b42
	13'h05a2: q2 = 16'h000a; // 0x0b44
	13'h05a3: q2 = 16'h200b; // 0x0b46
	13'h05a4: q2 = 16'h5080; // 0x0b48
	13'h05a5: q2 = 16'h2e80; // 0x0b4a
	13'h05a6: q2 = 16'h4eb9; // 0x0b4c
	13'h05a7: q2 = 16'h0000; // 0x0b4e
	13'h05a8: q2 = 16'h072e; // 0x0b50
	13'h05a9: q2 = 16'h3a00; // 0x0b52
	13'h05aa: q2 = 16'h4a79; // 0x0b54
	13'h05ab: q2 = 16'h0001; // 0x0b56
	13'h05ac: q2 = 16'h7fc6; // 0x0b58
	13'h05ad: q2 = 16'h6600; // 0x0b5a
	13'h05ae: q2 = 16'h0088; // 0x0b5c
	13'h05af: q2 = 16'h202c; // 0x0b5e
	13'h05b0: q2 = 16'h0004; // 0x0b60
	13'h05b1: q2 = 16'hb0b9; // 0x0b62
	13'h05b2: q2 = 16'h0001; // 0x0b64
	13'h05b3: q2 = 16'h7f64; // 0x0b66
	13'h05b4: q2 = 16'h6e0c; // 0x0b68
	13'h05b5: q2 = 16'h202b; // 0x0b6a
	13'h05b6: q2 = 16'h0004; // 0x0b6c
	13'h05b7: q2 = 16'hb0b9; // 0x0b6e
	13'h05b8: q2 = 16'h0001; // 0x0b70
	13'h05b9: q2 = 16'h7f64; // 0x0b72
	13'h05ba: q2 = 16'h6f6e; // 0x0b74
	13'h05bb: q2 = 16'h202c; // 0x0b76
	13'h05bc: q2 = 16'h0004; // 0x0b78
	13'h05bd: q2 = 16'hb0ab; // 0x0b7a
	13'h05be: q2 = 16'h0004; // 0x0b7c
	13'h05bf: q2 = 16'h6f32; // 0x0b7e
	13'h05c0: q2 = 16'h2ebc; // 0x0b80
	13'h05c1: q2 = 16'h0000; // 0x0b82
	13'h05c2: q2 = 16'hf80a; // 0x0b84
	13'h05c3: q2 = 16'h200e; // 0x0b86
	13'h05c4: q2 = 16'hd0bc; // 0x0b88
	13'h05c5: q2 = 16'hffff; // 0x0b8a
	13'h05c6: q2 = 16'hfff0; // 0x0b8c
	13'h05c7: q2 = 16'h2f00; // 0x0b8e
	13'h05c8: q2 = 16'h4eb9; // 0x0b90
	13'h05c9: q2 = 16'h0000; // 0x0b92
	13'h05ca: q2 = 16'h0750; // 0x0b94
	13'h05cb: q2 = 16'h4a9f; // 0x0b96
	13'h05cc: q2 = 16'h200c; // 0x0b98
	13'h05cd: q2 = 16'h5080; // 0x0b9a
	13'h05ce: q2 = 16'h2e80; // 0x0b9c
	13'h05cf: q2 = 16'h200e; // 0x0b9e
	13'h05d0: q2 = 16'hd0bc; // 0x0ba0
	13'h05d1: q2 = 16'hffff; // 0x0ba2
	13'h05d2: q2 = 16'hfff0; // 0x0ba4
	13'h05d3: q2 = 16'h2f00; // 0x0ba6
	13'h05d4: q2 = 16'h4eb9; // 0x0ba8
	13'h05d5: q2 = 16'h0000; // 0x0baa
	13'h05d6: q2 = 16'h0770; // 0x0bac
	13'h05d7: q2 = 16'h4a9f; // 0x0bae
	13'h05d8: q2 = 16'h6030; // 0x0bb0
	13'h05d9: q2 = 16'h2ebc; // 0x0bb2
	13'h05da: q2 = 16'h0000; // 0x0bb4
	13'h05db: q2 = 16'hf80f; // 0x0bb6
	13'h05dc: q2 = 16'h200e; // 0x0bb8
	13'h05dd: q2 = 16'hd0bc; // 0x0bba
	13'h05de: q2 = 16'hffff; // 0x0bbc
	13'h05df: q2 = 16'hfff0; // 0x0bbe
	13'h05e0: q2 = 16'h2f00; // 0x0bc0
	13'h05e1: q2 = 16'h4eb9; // 0x0bc2
	13'h05e2: q2 = 16'h0000; // 0x0bc4
	13'h05e3: q2 = 16'h0750; // 0x0bc6
	13'h05e4: q2 = 16'h4a9f; // 0x0bc8
	13'h05e5: q2 = 16'h200b; // 0x0bca
	13'h05e6: q2 = 16'h5080; // 0x0bcc
	13'h05e7: q2 = 16'h2e80; // 0x0bce
	13'h05e8: q2 = 16'h200e; // 0x0bd0
	13'h05e9: q2 = 16'hd0bc; // 0x0bd2
	13'h05ea: q2 = 16'hffff; // 0x0bd4
	13'h05eb: q2 = 16'hfff0; // 0x0bd6
	13'h05ec: q2 = 16'h2f00; // 0x0bd8
	13'h05ed: q2 = 16'h4eb9; // 0x0bda
	13'h05ee: q2 = 16'h0000; // 0x0bdc
	13'h05ef: q2 = 16'h0770; // 0x0bde
	13'h05f0: q2 = 16'h4a9f; // 0x0be0
	13'h05f1: q2 = 16'h6052; // 0x0be2
	13'h05f2: q2 = 16'h4247; // 0x0be4
	13'h05f3: q2 = 16'h4bee; // 0x0be6
	13'h05f4: q2 = 16'hfff0; // 0x0be8
	13'h05f5: q2 = 16'hbe7c; // 0x0bea
	13'h05f6: q2 = 16'h0003; // 0x0bec
	13'h05f7: q2 = 16'h6c14; // 0x0bee
	13'h05f8: q2 = 16'h3007; // 0x0bf0
	13'h05f9: q2 = 16'h48c0; // 0x0bf2
	13'h05fa: q2 = 16'hd0bc; // 0x0bf4
	13'h05fb: q2 = 16'h0001; // 0x0bf6
	13'h05fc: q2 = 16'h7ba8; // 0x0bf8
	13'h05fd: q2 = 16'h2040; // 0x0bfa
	13'h05fe: q2 = 16'h1a90; // 0x0bfc
	13'h05ff: q2 = 16'h5247; // 0x0bfe
	13'h0600: q2 = 16'h528d; // 0x0c00
	13'h0601: q2 = 16'h60e6; // 0x0c02
	13'h0602: q2 = 16'h4215; // 0x0c04
	13'h0603: q2 = 16'h2ebc; // 0x0c06
	13'h0604: q2 = 16'h0000; // 0x0c08
	13'h0605: q2 = 16'hf814; // 0x0c0a
	13'h0606: q2 = 16'h200e; // 0x0c0c
	13'h0607: q2 = 16'hd0bc; // 0x0c0e
	13'h0608: q2 = 16'hffff; // 0x0c10
	13'h0609: q2 = 16'hfff0; // 0x0c12
	13'h060a: q2 = 16'h2f00; // 0x0c14
	13'h060b: q2 = 16'h4eb9; // 0x0c16
	13'h060c: q2 = 16'h0000; // 0x0c18
	13'h060d: q2 = 16'h0770; // 0x0c1a
	13'h060e: q2 = 16'h4a9f; // 0x0c1c
	13'h060f: q2 = 16'h2ebc; // 0x0c1e
	13'h0610: q2 = 16'h0001; // 0x0c20
	13'h0611: q2 = 16'h860e; // 0x0c22
	13'h0612: q2 = 16'h200e; // 0x0c24
	13'h0613: q2 = 16'hd0bc; // 0x0c26
	13'h0614: q2 = 16'hffff; // 0x0c28
	13'h0615: q2 = 16'hfff0; // 0x0c2a
	13'h0616: q2 = 16'h2f00; // 0x0c2c
	13'h0617: q2 = 16'h4eb9; // 0x0c2e
	13'h0618: q2 = 16'h0000; // 0x0c30
	13'h0619: q2 = 16'h0770; // 0x0c32
	13'h061a: q2 = 16'h4a9f; // 0x0c34
	13'h061b: q2 = 16'h200e; // 0x0c36
	13'h061c: q2 = 16'hd0bc; // 0x0c38
	13'h061d: q2 = 16'hffff; // 0x0c3a
	13'h061e: q2 = 16'hfff0; // 0x0c3c
	13'h061f: q2 = 16'h2e80; // 0x0c3e
	13'h0620: q2 = 16'h4eb9; // 0x0c40
	13'h0621: q2 = 16'h0000; // 0x0c42
	13'h0622: q2 = 16'h072e; // 0x0c44
	13'h0623: q2 = 16'h3800; // 0x0c46
	13'h0624: q2 = 16'h3004; // 0x0c48
	13'h0625: q2 = 16'hd046; // 0x0c4a
	13'h0626: q2 = 16'hb07c; // 0x0c4c
	13'h0627: q2 = 16'h0016; // 0x0c4e
	13'h0628: q2 = 16'h6e0a; // 0x0c50
	13'h0629: q2 = 16'h3004; // 0x0c52
	13'h062a: q2 = 16'hd045; // 0x0c54
	13'h062b: q2 = 16'hb07c; // 0x0c56
	13'h062c: q2 = 16'h0016; // 0x0c58
	13'h062d: q2 = 16'h6f1c; // 0x0c5a
	13'h062e: q2 = 16'h200e; // 0x0c5c
	13'h062f: q2 = 16'hd0bc; // 0x0c5e
	13'h0630: q2 = 16'hffff; // 0x0c60
	13'h0631: q2 = 16'hfff4; // 0x0c62
	13'h0632: q2 = 16'h2e80; // 0x0c64
	13'h0633: q2 = 16'h200e; // 0x0c66
	13'h0634: q2 = 16'hd0bc; // 0x0c68
	13'h0635: q2 = 16'hffff; // 0x0c6a
	13'h0636: q2 = 16'hfff0; // 0x0c6c
	13'h0637: q2 = 16'h2f00; // 0x0c6e
	13'h0638: q2 = 16'h4eb9; // 0x0c70
	13'h0639: q2 = 16'h0000; // 0x0c72
	13'h063a: q2 = 16'h0750; // 0x0c74
	13'h063b: q2 = 16'h4a9f; // 0x0c76
	13'h063c: q2 = 16'h3ebc; // 0x0c78
	13'h063d: q2 = 16'h0026; // 0x0c7a
	13'h063e: q2 = 16'h4267; // 0x0c7c
	13'h063f: q2 = 16'h3f3c; // 0x0c7e
	13'h0640: q2 = 16'h0064; // 0x0c80
	13'h0641: q2 = 16'h3f3c; // 0x0c82
	13'h0642: q2 = 16'h001f; // 0x0c84
	13'h0643: q2 = 16'h200e; // 0x0c86
	13'h0644: q2 = 16'hd0bc; // 0x0c88
	13'h0645: q2 = 16'hffff; // 0x0c8a
	13'h0646: q2 = 16'hfff0; // 0x0c8c
	13'h0647: q2 = 16'h2f00; // 0x0c8e
	13'h0648: q2 = 16'h4eb9; // 0x0c90
	13'h0649: q2 = 16'h0000; // 0x0c92
	13'h064a: q2 = 16'h026c; // 0x0c94
	13'h064b: q2 = 16'hdefc; // 0x0c96
	13'h064c: q2 = 16'h000a; // 0x0c98
	13'h064d: q2 = 16'h4a9f; // 0x0c9a
	13'h064e: q2 = 16'h4cdf; // 0x0c9c
	13'h064f: q2 = 16'h38f0; // 0x0c9e
	13'h0650: q2 = 16'h4e5e; // 0x0ca0
	13'h0651: q2 = 16'h4e75; // 0x0ca2
	13'h0652: q2 = 16'h4e56; // 0x0ca4
	13'h0653: q2 = 16'h0000; // 0x0ca6
	13'h0654: q2 = 16'h48e7; // 0x0ca8
	13'h0655: q2 = 16'h0704; // 0x0caa
	13'h0656: q2 = 16'h2a79; // 0x0cac
	13'h0657: q2 = 16'h0001; // 0x0cae
	13'h0658: q2 = 16'h7fb8; // 0x0cb0
	13'h0659: q2 = 16'h0c55; // 0x0cb2
	13'h065a: q2 = 16'h0003; // 0x0cb4
	13'h065b: q2 = 16'h6e08; // 0x0cb6
	13'h065c: q2 = 16'h33fc; // 0x0cb8
	13'h065d: q2 = 16'h7d0e; // 0x0cba
	13'h065e: q2 = 16'h0001; // 0x0cbc
	13'h065f: q2 = 16'h8a76; // 0x0cbe
	13'h0660: q2 = 16'h33f9; // 0x0cc0
	13'h0661: q2 = 16'h0001; // 0x0cc2
	13'h0662: q2 = 16'h8a76; // 0x0cc4
	13'h0663: q2 = 16'h0001; // 0x0cc6
	13'h0664: q2 = 16'h7eba; // 0x0cc8
	13'h0665: q2 = 16'h4eb9; // 0x0cca
	13'h0666: q2 = 16'h0000; // 0x0ccc
	13'h0667: q2 = 16'h0226; // 0x0cce
	13'h0668: q2 = 16'h4eb9; // 0x0cd0
	13'h0669: q2 = 16'h0000; // 0x0cd2
	13'h066a: q2 = 16'h0ea2; // 0x0cd4
	13'h066b: q2 = 16'h4eb9; // 0x0cd6
	13'h066c: q2 = 16'h0000; // 0x0cd8
	13'h066d: q2 = 16'h41ae; // 0x0cda
	13'h066e: q2 = 16'h4eb9; // 0x0cdc
	13'h066f: q2 = 16'h0000; // 0x0cde
	13'h0670: q2 = 16'hb3c6; // 0x0ce0
	13'h0671: q2 = 16'h4eb9; // 0x0ce2
	13'h0672: q2 = 16'h0000; // 0x0ce4
	13'h0673: q2 = 16'h1e8a; // 0x0ce6
	13'h0674: q2 = 16'h4eb9; // 0x0ce8
	13'h0675: q2 = 16'h0000; // 0x0cea
	13'h0676: q2 = 16'h4dee; // 0x0cec
	13'h0677: q2 = 16'h4a79; // 0x0cee
	13'h0678: q2 = 16'h0001; // 0x0cf0
	13'h0679: q2 = 16'h7fc8; // 0x0cf2
	13'h067a: q2 = 16'h670e; // 0x0cf4
	13'h067b: q2 = 16'h3eb9; // 0x0cf6
	13'h067c: q2 = 16'h0001; // 0x0cf8
	13'h067d: q2 = 16'h8054; // 0x0cfa
	13'h067e: q2 = 16'h5257; // 0x0cfc
	13'h067f: q2 = 16'h4eb9; // 0x0cfe
	13'h0680: q2 = 16'h0000; // 0x0d00
	13'h0681: q2 = 16'h8856; // 0x0d02
	13'h0682: q2 = 16'h4279; // 0x0d04
	13'h0683: q2 = 16'h0001; // 0x0d06
	13'h0684: q2 = 16'h7fc8; // 0x0d08
	13'h0685: q2 = 16'h4eb9; // 0x0d0a
	13'h0686: q2 = 16'h0000; // 0x0d0c
	13'h0687: q2 = 16'h8330; // 0x0d0e
	13'h0688: q2 = 16'h4eb9; // 0x0d10
	13'h0689: q2 = 16'h0000; // 0x0d12
	13'h068a: q2 = 16'h5a9c; // 0x0d14
	13'h068b: q2 = 16'h4eb9; // 0x0d16
	13'h068c: q2 = 16'h0000; // 0x0d18
	13'h068d: q2 = 16'h2cba; // 0x0d1a
	13'h068e: q2 = 16'h4a79; // 0x0d1c
	13'h068f: q2 = 16'h0001; // 0x0d1e
	13'h0690: q2 = 16'h7eb8; // 0x0d20
	13'h0691: q2 = 16'h670e; // 0x0d22
	13'h0692: q2 = 16'h2ebc; // 0x0d24
	13'h0693: q2 = 16'h0000; // 0x0d26
	13'h0694: q2 = 16'hf376; // 0x0d28
	13'h0695: q2 = 16'h4eb9; // 0x0d2a
	13'h0696: q2 = 16'h0000; // 0x0d2c
	13'h0697: q2 = 16'h7ff8; // 0x0d2e
	13'h0698: q2 = 16'h600c; // 0x0d30
	13'h0699: q2 = 16'h2ebc; // 0x0d32
	13'h069a: q2 = 16'h0000; // 0x0d34
	13'h069b: q2 = 16'hfaf6; // 0x0d36
	13'h069c: q2 = 16'h4eb9; // 0x0d38
	13'h069d: q2 = 16'h0000; // 0x0d3a
	13'h069e: q2 = 16'h7ff8; // 0x0d3c
	13'h069f: q2 = 16'h4279; // 0x0d3e
	13'h06a0: q2 = 16'h0001; // 0x0d40
	13'h06a1: q2 = 16'h7eb8; // 0x0d42
	13'h06a2: q2 = 16'h4eb9; // 0x0d44
	13'h06a3: q2 = 16'h0000; // 0x0d46
	13'h06a4: q2 = 16'h90d4; // 0x0d48
	13'h06a5: q2 = 16'h33fc; // 0x0d4a
	13'h06a6: q2 = 16'h0001; // 0x0d4c
	13'h06a7: q2 = 16'h0001; // 0x0d4e
	13'h06a8: q2 = 16'h7b9e; // 0x0d50
	13'h06a9: q2 = 16'h7e3c; // 0x0d52
	13'h06aa: q2 = 16'h4a47; // 0x0d54
	13'h06ab: q2 = 16'h6724; // 0x0d56
	13'h06ac: q2 = 16'h23fc; // 0x0d58
	13'h06ad: q2 = 16'h0000; // 0x0d5a
	13'h06ae: q2 = 16'h0002; // 0x0d5c
	13'h06af: q2 = 16'h0001; // 0x0d5e
	13'h06b0: q2 = 16'h7fc2; // 0x0d60
	13'h06b1: q2 = 16'h4eb9; // 0x0d62
	13'h06b2: q2 = 16'h0000; // 0x0d64
	13'h06b3: q2 = 16'h4820; // 0x0d66
	13'h06b4: q2 = 16'h4eb9; // 0x0d68
	13'h06b5: q2 = 16'h0000; // 0x0d6a
	13'h06b6: q2 = 16'h18d0; // 0x0d6c
	13'h06b7: q2 = 16'h4ab9; // 0x0d6e
	13'h06b8: q2 = 16'h0001; // 0x0d70
	13'h06b9: q2 = 16'h7fc2; // 0x0d72
	13'h06ba: q2 = 16'h6702; // 0x0d74
	13'h06bb: q2 = 16'h60f6; // 0x0d76
	13'h06bc: q2 = 16'h5347; // 0x0d78
	13'h06bd: q2 = 16'h60d8; // 0x0d7a
	13'h06be: q2 = 16'h4279; // 0x0d7c
	13'h06bf: q2 = 16'h0001; // 0x0d7e
	13'h06c0: q2 = 16'h7b9e; // 0x0d80
	13'h06c1: q2 = 16'h23fc; // 0x0d82
	13'h06c2: q2 = 16'h0000; // 0x0d84
	13'h06c3: q2 = 16'h0002; // 0x0d86
	13'h06c4: q2 = 16'h0001; // 0x0d88
	13'h06c5: q2 = 16'h7fc2; // 0x0d8a
	13'h06c6: q2 = 16'h33fc; // 0x0d8c
	13'h06c7: q2 = 16'h0001; // 0x0d8e
	13'h06c8: q2 = 16'h0001; // 0x0d90
	13'h06c9: q2 = 16'h805a; // 0x0d92
	13'h06ca: q2 = 16'h4eb9; // 0x0d94
	13'h06cb: q2 = 16'h0000; // 0x0d96
	13'h06cc: q2 = 16'h3434; // 0x0d98
	13'h06cd: q2 = 16'h4eb9; // 0x0d9a
	13'h06ce: q2 = 16'h0000; // 0x0d9c
	13'h06cf: q2 = 16'h18d0; // 0x0d9e
	13'h06d0: q2 = 16'h4eb9; // 0x0da0
	13'h06d1: q2 = 16'h0000; // 0x0da2
	13'h06d2: q2 = 16'h4820; // 0x0da4
	13'h06d3: q2 = 16'h4eb9; // 0x0da6
	13'h06d4: q2 = 16'h0000; // 0x0da8
	13'h06d5: q2 = 16'h909e; // 0x0daa
	13'h06d6: q2 = 16'h4eb9; // 0x0dac
	13'h06d7: q2 = 16'h0000; // 0x0dae
	13'h06d8: q2 = 16'h3fcc; // 0x0db0
	13'h06d9: q2 = 16'h4eb9; // 0x0db2
	13'h06da: q2 = 16'h0000; // 0x0db4
	13'h06db: q2 = 16'h3396; // 0x0db6
	13'h06dc: q2 = 16'h4a40; // 0x0db8
	13'h06dd: q2 = 16'h6726; // 0x0dba
	13'h06de: q2 = 16'h4eb9; // 0x0dbc
	13'h06df: q2 = 16'h0000; // 0x0dbe
	13'h06e0: q2 = 16'h4738; // 0x0dc0
	13'h06e1: q2 = 16'h4a40; // 0x0dc2
	13'h06e2: q2 = 16'h671c; // 0x0dc4
	13'h06e3: q2 = 16'h4eb9; // 0x0dc6
	13'h06e4: q2 = 16'h0000; // 0x0dc8
	13'h06e5: q2 = 16'h16c2; // 0x0dca
	13'h06e6: q2 = 16'h4a40; // 0x0dcc
	13'h06e7: q2 = 16'h6712; // 0x0dce
	13'h06e8: q2 = 16'h4eb9; // 0x0dd0
	13'h06e9: q2 = 16'h0000; // 0x0dd2
	13'h06ea: q2 = 16'h3fac; // 0x0dd4
	13'h06eb: q2 = 16'h4a40; // 0x0dd6
	13'h06ec: q2 = 16'h6708; // 0x0dd8
	13'h06ed: q2 = 16'h4eb9; // 0x0dda
	13'h06ee: q2 = 16'h0000; // 0x0ddc
	13'h06ef: q2 = 16'h18d0; // 0x0dde
	13'h06f0: q2 = 16'h600c; // 0x0de0
	13'h06f1: q2 = 16'h4ab9; // 0x0de2
	13'h06f2: q2 = 16'h0001; // 0x0de4
	13'h06f3: q2 = 16'h7fc2; // 0x0de6
	13'h06f4: q2 = 16'h6702; // 0x0de8
	13'h06f5: q2 = 16'h60f6; // 0x0dea
	13'h06f6: q2 = 16'h6094; // 0x0dec
	13'h06f7: q2 = 16'h4eb9; // 0x0dee
	13'h06f8: q2 = 16'h0000; // 0x0df0
	13'h06f9: q2 = 16'h4738; // 0x0df2
	13'h06fa: q2 = 16'hb07c; // 0x0df4
	13'h06fb: q2 = 16'h0001; // 0x0df6
	13'h06fc: q2 = 16'h6614; // 0x0df8
	13'h06fd: q2 = 16'h4eb9; // 0x0dfa
	13'h06fe: q2 = 16'h0000; // 0x0dfc
	13'h06ff: q2 = 16'h4ec6; // 0x0dfe
	13'h0700: q2 = 16'hb07c; // 0x0e00
	13'h0701: q2 = 16'h0001; // 0x0e02
	13'h0702: q2 = 16'h675c; // 0x0e04
	13'h0703: q2 = 16'h4eb9; // 0x0e06
	13'h0704: q2 = 16'h0000; // 0x0e08
	13'h0705: q2 = 16'ha792; // 0x0e0a
	13'h0706: q2 = 16'h6054; // 0x0e0c
	13'h0707: q2 = 16'h2eb9; // 0x0e0e
	13'h0708: q2 = 16'h0000; // 0x0e10
	13'h0709: q2 = 16'hf816; // 0x0e12
	13'h070a: q2 = 16'h4eb9; // 0x0e14
	13'h070b: q2 = 16'h0000; // 0x0e16
	13'h070c: q2 = 16'h3da4; // 0x0e18
	13'h070d: q2 = 16'h4eb9; // 0x0e1a
	13'h070e: q2 = 16'h0000; // 0x0e1c
	13'h070f: q2 = 16'h4446; // 0x0e1e
	13'h0710: q2 = 16'h3c15; // 0x0e20
	13'h0711: q2 = 16'he546; // 0x0e22
	13'h0712: q2 = 16'hdc55; // 0x0e24
	13'h0713: q2 = 16'hbc7c; // 0x0e26
	13'h0714: q2 = 16'h00fa; // 0x0e28
	13'h0715: q2 = 16'h6f04; // 0x0e2a
	13'h0716: q2 = 16'h3c3c; // 0x0e2c
	13'h0717: q2 = 16'h00fa; // 0x0e2e
	13'h0718: q2 = 16'h3e86; // 0x0e30
	13'h0719: q2 = 16'h4eb9; // 0x0e32
	13'h071a: q2 = 16'h0000; // 0x0e34
	13'h071b: q2 = 16'h8ee8; // 0x0e36
	13'h071c: q2 = 16'h4eb9; // 0x0e38
	13'h071d: q2 = 16'h0000; // 0x0e3a
	13'h071e: q2 = 16'h0db8; // 0x0e3c
	13'h071f: q2 = 16'h4eb9; // 0x0e3e
	13'h0720: q2 = 16'h0000; // 0x0e40
	13'h0721: q2 = 16'h6b28; // 0x0e42
	13'h0722: q2 = 16'h3b7c; // 0x0e44
	13'h0723: q2 = 16'hffff; // 0x0e46
	13'h0724: q2 = 16'h0024; // 0x0e48
	13'h0725: q2 = 16'h0c55; // 0x0e4a
	13'h0726: q2 = 16'h007d; // 0x0e4c
	13'h0727: q2 = 16'h6c02; // 0x0e4e
	13'h0728: q2 = 16'h5255; // 0x0e50
	13'h0729: q2 = 16'h2eb9; // 0x0e52
	13'h072a: q2 = 16'h0000; // 0x0e54
	13'h072b: q2 = 16'hf81a; // 0x0e56
	13'h072c: q2 = 16'h4eb9; // 0x0e58
	13'h072d: q2 = 16'h0000; // 0x0e5a
	13'h072e: q2 = 16'h3da4; // 0x0e5c
	13'h072f: q2 = 16'h6000; // 0x0e5e
	13'h0730: q2 = 16'hfe52; // 0x0e60
	13'h0731: q2 = 16'h4a9f; // 0x0e62
	13'h0732: q2 = 16'h4cdf; // 0x0e64
	13'h0733: q2 = 16'h20c0; // 0x0e66
	13'h0734: q2 = 16'h4e5e; // 0x0e68
	13'h0735: q2 = 16'h4e75; // 0x0e6a
	13'h0736: q2 = 16'h4e56; // 0x0e6c
	13'h0737: q2 = 16'hfffc; // 0x0e6e
	13'h0738: q2 = 16'h4280; // 0x0e70
	13'h0739: q2 = 16'h3039; // 0x0e72
	13'h073a: q2 = 16'h0001; // 0x0e74
	13'h073b: q2 = 16'h8a76; // 0x0e76
	13'h073c: q2 = 16'hc0fc; // 0x0e78
	13'h073d: q2 = 16'h873d; // 0x0e7a
	13'h073e: q2 = 16'hd0bc; // 0x0e7c
	13'h073f: q2 = 16'h0000; // 0x0e7e
	13'h0740: q2 = 16'h3619; // 0x0e80
	13'h0741: q2 = 16'h33c0; // 0x0e82
	13'h0742: q2 = 16'h0001; // 0x0e84
	13'h0743: q2 = 16'h8a76; // 0x0e86
	13'h0744: q2 = 16'h4280; // 0x0e88
	13'h0745: q2 = 16'h302e; // 0x0e8a
	13'h0746: q2 = 16'h000a; // 0x0e8c
	13'h0747: q2 = 16'h906e; // 0x0e8e
	13'h0748: q2 = 16'h0008; // 0x0e90
	13'h0749: q2 = 16'h5240; // 0x0e92
	13'h074a: q2 = 16'hc0f9; // 0x0e94
	13'h074b: q2 = 16'h0001; // 0x0e96
	13'h074c: q2 = 16'h8a76; // 0x0e98
	13'h074d: q2 = 16'h4281; // 0x0e9a
	13'h074e: q2 = 16'h7210; // 0x0e9c
	13'h074f: q2 = 16'he2a8; // 0x0e9e
	13'h0750: q2 = 16'hd06e; // 0x0ea0
	13'h0751: q2 = 16'h0008; // 0x0ea2
	13'h0752: q2 = 16'h4e5e; // 0x0ea4
	13'h0753: q2 = 16'h4e75; // 0x0ea6
	13'h0754: q2 = 16'h4e56; // 0x0ea8
	13'h0755: q2 = 16'h0000; // 0x0eaa
	13'h0756: q2 = 16'h48e7; // 0x0eac
	13'h0757: q2 = 16'h030c; // 0x0eae
	13'h0758: q2 = 16'h287c; // 0x0eb0
	13'h0759: q2 = 16'h0000; // 0x0eb2
	13'h075a: q2 = 16'hf81e; // 0x0eb4
	13'h075b: q2 = 16'h2a7c; // 0x0eb6
	13'h075c: q2 = 16'h0001; // 0x0eb8
	13'h075d: q2 = 16'h75e8; // 0x0eba
	13'h075e: q2 = 16'h4247; // 0x0ebc
	13'h075f: q2 = 16'hbe7c; // 0x0ebe
	13'h0760: q2 = 16'h0100; // 0x0ec0
	13'h0761: q2 = 16'h6c1a; // 0x0ec2
	13'h0762: q2 = 16'h3007; // 0x0ec4
	13'h0763: q2 = 16'hc07c; // 0x0ec6
	13'h0764: q2 = 16'h0003; // 0x0ec8
	13'h0765: q2 = 16'h6604; // 0x0eca
	13'h0766: q2 = 16'h4255; // 0x0ecc
	13'h0767: q2 = 16'h6008; // 0x0ece
	13'h0768: q2 = 16'h1014; // 0x0ed0
	13'h0769: q2 = 16'h4880; // 0x0ed2
	13'h076a: q2 = 16'h3a80; // 0x0ed4
	13'h076b: q2 = 16'h528c; // 0x0ed6
	13'h076c: q2 = 16'h5247; // 0x0ed8
	13'h076d: q2 = 16'h548d; // 0x0eda
	13'h076e: q2 = 16'h60e0; // 0x0edc
	13'h076f: q2 = 16'h4a9f; // 0x0ede
	13'h0770: q2 = 16'h4cdf; // 0x0ee0
	13'h0771: q2 = 16'h3080; // 0x0ee2
	13'h0772: q2 = 16'h4e5e; // 0x0ee4
	13'h0773: q2 = 16'h4e75; // 0x0ee6
	13'h0774: q2 = 16'h4e56; // 0x0ee8
	13'h0775: q2 = 16'hfff4; // 0x0eea
	13'h0776: q2 = 16'h48e7; // 0x0eec
	13'h0777: q2 = 16'h0104; // 0x0eee
	13'h0778: q2 = 16'h4a79; // 0x0ef0
	13'h0779: q2 = 16'h0001; // 0x0ef2
	13'h077a: q2 = 16'h7fc6; // 0x0ef4
	13'h077b: q2 = 16'h6600; // 0x0ef6
	13'h077c: q2 = 16'h017a; // 0x0ef8
	13'h077d: q2 = 16'h4a79; // 0x0efa
	13'h077e: q2 = 16'h0001; // 0x0efc
	13'h077f: q2 = 16'h8676; // 0x0efe
	13'h0780: q2 = 16'h6600; // 0x0f00
	13'h0781: q2 = 16'h0170; // 0x0f02
	13'h0782: q2 = 16'h4a79; // 0x0f04
	13'h0783: q2 = 16'h0001; // 0x0f06
	13'h0784: q2 = 16'h7faa; // 0x0f08
	13'h0785: q2 = 16'h6600; // 0x0f0a
	13'h0786: q2 = 16'h0166; // 0x0f0c
	13'h0787: q2 = 16'h2a79; // 0x0f0e
	13'h0788: q2 = 16'h0001; // 0x0f10
	13'h0789: q2 = 16'h7fb8; // 0x0f12
	13'h078a: q2 = 16'h200e; // 0x0f14
	13'h078b: q2 = 16'hd0bc; // 0x0f16
	13'h078c: q2 = 16'hffff; // 0x0f18
	13'h078d: q2 = 16'hfff4; // 0x0f1a
	13'h078e: q2 = 16'h2e80; // 0x0f1c
	13'h078f: q2 = 16'h3f2e; // 0x0f1e
	13'h0790: q2 = 16'h0008; // 0x0f20
	13'h0791: q2 = 16'h4eb9; // 0x0f22
	13'h0792: q2 = 16'h0000; // 0x0f24
	13'h0793: q2 = 16'h0828; // 0x0f26
	13'h0794: q2 = 16'h4a5f; // 0x0f28
	13'h0795: q2 = 16'h2ebc; // 0x0f2a
	13'h0796: q2 = 16'h0000; // 0x0f2c
	13'h0797: q2 = 16'hf8e6; // 0x0f2e
	13'h0798: q2 = 16'h200e; // 0x0f30
	13'h0799: q2 = 16'hd0bc; // 0x0f32
	13'h079a: q2 = 16'hffff; // 0x0f34
	13'h079b: q2 = 16'hfff4; // 0x0f36
	13'h079c: q2 = 16'h2f00; // 0x0f38
	13'h079d: q2 = 16'h4eb9; // 0x0f3a
	13'h079e: q2 = 16'h0000; // 0x0f3c
	13'h079f: q2 = 16'h0770; // 0x0f3e
	13'h07a0: q2 = 16'h4a9f; // 0x0f40
	13'h07a1: q2 = 16'h4aad; // 0x0f42
	13'h07a2: q2 = 16'h0004; // 0x0f44
	13'h07a3: q2 = 16'h671a; // 0x0f46
	13'h07a4: q2 = 16'h200e; // 0x0f48
	13'h07a5: q2 = 16'hd0bc; // 0x0f4a
	13'h07a6: q2 = 16'hffff; // 0x0f4c
	13'h07a7: q2 = 16'hfff4; // 0x0f4e
	13'h07a8: q2 = 16'h2e80; // 0x0f50
	13'h07a9: q2 = 16'h200d; // 0x0f52
	13'h07aa: q2 = 16'h5080; // 0x0f54
	13'h07ab: q2 = 16'h2f00; // 0x0f56
	13'h07ac: q2 = 16'h4eb9; // 0x0f58
	13'h07ad: q2 = 16'h0000; // 0x0f5a
	13'h07ae: q2 = 16'h0908; // 0x0f5c
	13'h07af: q2 = 16'h4a9f; // 0x0f5e
	13'h07b0: q2 = 16'h6018; // 0x0f60
	13'h07b1: q2 = 16'h200e; // 0x0f62
	13'h07b2: q2 = 16'hd0bc; // 0x0f64
	13'h07b3: q2 = 16'hffff; // 0x0f66
	13'h07b4: q2 = 16'hfff4; // 0x0f68
	13'h07b5: q2 = 16'h2e80; // 0x0f6a
	13'h07b6: q2 = 16'h200d; // 0x0f6c
	13'h07b7: q2 = 16'h5080; // 0x0f6e
	13'h07b8: q2 = 16'h2f00; // 0x0f70
	13'h07b9: q2 = 16'h4eb9; // 0x0f72
	13'h07ba: q2 = 16'h0000; // 0x0f74
	13'h07bb: q2 = 16'h0750; // 0x0f76
	13'h07bc: q2 = 16'h4a9f; // 0x0f78
	13'h07bd: q2 = 16'h302e; // 0x0f7a
	13'h07be: q2 = 16'h0008; // 0x0f7c
	13'h07bf: q2 = 16'h48c0; // 0x0f7e
	13'h07c0: q2 = 16'hd1ad; // 0x0f80
	13'h07c1: q2 = 16'h0004; // 0x0f82
	13'h07c2: q2 = 16'h2039; // 0x0f84
	13'h07c3: q2 = 16'h0000; // 0x0f86
	13'h07c4: q2 = 16'hf8de; // 0x0f88
	13'h07c5: q2 = 16'hb0ad; // 0x0f8a
	13'h07c6: q2 = 16'h0004; // 0x0f8c
	13'h07c7: q2 = 16'h6c5e; // 0x0f8e
	13'h07c8: q2 = 16'h2039; // 0x0f90
	13'h07c9: q2 = 16'h0000; // 0x0f92
	13'h07ca: q2 = 16'hf8e2; // 0x0f94
	13'h07cb: q2 = 16'h91ad; // 0x0f96
	13'h07cc: q2 = 16'h0004; // 0x0f98
	13'h07cd: q2 = 16'h200d; // 0x0f9a
	13'h07ce: q2 = 16'h5080; // 0x0f9c
	13'h07cf: q2 = 16'h2e80; // 0x0f9e
	13'h07d0: q2 = 16'h2f2d; // 0x0fa0
	13'h07d1: q2 = 16'h0004; // 0x0fa2
	13'h07d2: q2 = 16'h4eb9; // 0x0fa4
	13'h07d3: q2 = 16'h0000; // 0x0fa6
	13'h07d4: q2 = 16'h0892; // 0x0fa8
	13'h07d5: q2 = 16'h4a9f; // 0x0faa
	13'h07d6: q2 = 16'h2ebc; // 0x0fac
	13'h07d7: q2 = 16'h0000; // 0x0fae
	13'h07d8: q2 = 16'hf8e9; // 0x0fb0
	13'h07d9: q2 = 16'h200d; // 0x0fb2
	13'h07da: q2 = 16'h5080; // 0x0fb4
	13'h07db: q2 = 16'h2f00; // 0x0fb6
	13'h07dc: q2 = 16'h4eb9; // 0x0fb8
	13'h07dd: q2 = 16'h0000; // 0x0fba
	13'h07de: q2 = 16'h0770; // 0x0fbc
	13'h07df: q2 = 16'h4a9f; // 0x0fbe
	13'h07e0: q2 = 16'h3ebc; // 0x0fc0
	13'h07e1: q2 = 16'h001f; // 0x0fc2
	13'h07e2: q2 = 16'h3f3c; // 0x0fc4
	13'h07e3: q2 = 16'h001f; // 0x0fc6
	13'h07e4: q2 = 16'h4eb9; // 0x0fc8
	13'h07e5: q2 = 16'h0000; // 0x0fca
	13'h07e6: q2 = 16'h01e4; // 0x0fcc
	13'h07e7: q2 = 16'h4a5f; // 0x0fce
	13'h07e8: q2 = 16'h4a79; // 0x0fd0
	13'h07e9: q2 = 16'h0001; // 0x0fd2
	13'h07ea: q2 = 16'h7582; // 0x0fd4
	13'h07eb: q2 = 16'h6f16; // 0x0fd6
	13'h07ec: q2 = 16'h4eb9; // 0x0fd8
	13'h07ed: q2 = 16'h0000; // 0x0fda
	13'h07ee: q2 = 16'h0d7c; // 0x0fdc
	13'h07ef: q2 = 16'h52b9; // 0x0fde
	13'h07f0: q2 = 16'h0001; // 0x0fe0
	13'h07f1: q2 = 16'h75b6; // 0x0fe2
	13'h07f2: q2 = 16'h3079; // 0x0fe4
	13'h07f3: q2 = 16'h0001; // 0x0fe6
	13'h07f4: q2 = 16'h7582; // 0x0fe8
	13'h07f5: q2 = 16'h2b48; // 0x0fea
	13'h07f6: q2 = 16'h0018; // 0x0fec
	13'h07f7: q2 = 16'h3079; // 0x0fee
	13'h07f8: q2 = 16'h0001; // 0x0ff0
	13'h07f9: q2 = 16'h7580; // 0x0ff2
	13'h07fa: q2 = 16'hb1ed; // 0x0ff4
	13'h07fb: q2 = 16'h0018; // 0x0ff6
	13'h07fc: q2 = 16'h6646; // 0x0ff8
	13'h07fd: q2 = 16'h3079; // 0x0ffa
	13'h07fe: q2 = 16'h0001; // 0x0ffc
	13'h07ff: q2 = 16'h7580; // 0x0ffe
	13'h0800: q2 = 16'hb1ed; // 0x1000
	13'h0801: q2 = 16'h0004; // 0x1002
	13'h0802: q2 = 16'h6e3a; // 0x1004
	13'h0803: q2 = 16'h4a79; // 0x1006
	13'h0804: q2 = 16'h0001; // 0x1008
	13'h0805: q2 = 16'h7580; // 0x100a
	13'h0806: q2 = 16'h6f32; // 0x100c
	13'h0807: q2 = 16'h4eb9; // 0x100e
	13'h0808: q2 = 16'h0000; // 0x1010
	13'h0809: q2 = 16'h0d7c; // 0x1012
	13'h080a: q2 = 16'h52b9; // 0x1014
	13'h080b: q2 = 16'h0001; // 0x1016
	13'h080c: q2 = 16'h75b2; // 0x1018
	13'h080d: q2 = 16'h3039; // 0x101a
	13'h080e: q2 = 16'h0001; // 0x101c
	13'h080f: q2 = 16'h7580; // 0x101e
	13'h0810: q2 = 16'hb079; // 0x1020
	13'h0811: q2 = 16'h0001; // 0x1022
	13'h0812: q2 = 16'h7582; // 0x1024
	13'h0813: q2 = 16'h660e; // 0x1026
	13'h0814: q2 = 16'h3039; // 0x1028
	13'h0815: q2 = 16'h0001; // 0x102a
	13'h0816: q2 = 16'h7582; // 0x102c
	13'h0817: q2 = 16'h48c0; // 0x102e
	13'h0818: q2 = 16'hd1ad; // 0x1030
	13'h0819: q2 = 16'h0018; // 0x1032
	13'h081a: q2 = 16'h600a; // 0x1034
	13'h081b: q2 = 16'h3079; // 0x1036
	13'h081c: q2 = 16'h0001; // 0x1038
	13'h081d: q2 = 16'h7582; // 0x103a
	13'h081e: q2 = 16'h2b48; // 0x103c
	13'h081f: q2 = 16'h0018; // 0x103e
	13'h0820: q2 = 16'h4a79; // 0x1040
	13'h0821: q2 = 16'h0001; // 0x1042
	13'h0822: q2 = 16'h7582; // 0x1044
	13'h0823: q2 = 16'h6f24; // 0x1046
	13'h0824: q2 = 16'h202d; // 0x1048
	13'h0825: q2 = 16'h0004; // 0x104a
	13'h0826: q2 = 16'hb0ad; // 0x104c
	13'h0827: q2 = 16'h0018; // 0x104e
	13'h0828: q2 = 16'h6d1a; // 0x1050
	13'h0829: q2 = 16'h4eb9; // 0x1052
	13'h082a: q2 = 16'h0000; // 0x1054
	13'h082b: q2 = 16'h0d7c; // 0x1056
	13'h082c: q2 = 16'h52b9; // 0x1058
	13'h082d: q2 = 16'h0001; // 0x105a
	13'h082e: q2 = 16'h75b6; // 0x105c
	13'h082f: q2 = 16'h3039; // 0x105e
	13'h0830: q2 = 16'h0001; // 0x1060
	13'h0831: q2 = 16'h7582; // 0x1062
	13'h0832: q2 = 16'h48c0; // 0x1064
	13'h0833: q2 = 16'hd1ad; // 0x1066
	13'h0834: q2 = 16'h0018; // 0x1068
	13'h0835: q2 = 16'h60dc; // 0x106a
	13'h0836: q2 = 16'h4eb9; // 0x106c
	13'h0837: q2 = 16'h0000; // 0x106e
	13'h0838: q2 = 16'h8a92; // 0x1070
	13'h0839: q2 = 16'h4a9f; // 0x1072
	13'h083a: q2 = 16'h4cdf; // 0x1074
	13'h083b: q2 = 16'h2000; // 0x1076
	13'h083c: q2 = 16'h4e5e; // 0x1078
	13'h083d: q2 = 16'h4e75; // 0x107a
	13'h083e: q2 = 16'h4e56; // 0x107c
	13'h083f: q2 = 16'hfffc; // 0x107e
	13'h0840: q2 = 16'h4a79; // 0x1080
	13'h0841: q2 = 16'h0001; // 0x1082
	13'h0842: q2 = 16'h8676; // 0x1084
	13'h0843: q2 = 16'h6704; // 0x1086
	13'h0844: q2 = 16'h4240; // 0x1088
	13'h0845: q2 = 16'h600e; // 0x108a
	13'h0846: q2 = 16'h4a79; // 0x108c
	13'h0847: q2 = 16'h0001; // 0x108e
	13'h0848: q2 = 16'h81fc; // 0x1090
	13'h0849: q2 = 16'h6604; // 0x1092
	13'h084a: q2 = 16'h7001; // 0x1094
	13'h084b: q2 = 16'h6002; // 0x1096
	13'h084c: q2 = 16'h4240; // 0x1098
	13'h084d: q2 = 16'h4e5e; // 0x109a
	13'h084e: q2 = 16'h4e75; // 0x109c
	13'h084f: q2 = 16'h4e56; // 0x109e
	13'h0850: q2 = 16'hfffc; // 0x10a0
	13'h0851: q2 = 16'h4ab9; // 0x10a2
	13'h0852: q2 = 16'h0001; // 0x10a4
	13'h0853: q2 = 16'h7fa2; // 0x10a6
	13'h0854: q2 = 16'h6626; // 0x10a8
	13'h0855: q2 = 16'h23f9; // 0x10aa
	13'h0856: q2 = 16'h0000; // 0x10ac
	13'h0857: q2 = 16'hf8ec; // 0x10ae
	13'h0858: q2 = 16'h0001; // 0x10b0
	13'h0859: q2 = 16'h7fa2; // 0x10b2
	13'h085a: q2 = 16'h4eb9; // 0x10b4
	13'h085b: q2 = 16'h0000; // 0x10b6
	13'h085c: q2 = 16'h907c; // 0x10b8
	13'h085d: q2 = 16'h4a40; // 0x10ba
	13'h085e: q2 = 16'h6612; // 0x10bc
	13'h085f: q2 = 16'h3039; // 0x10be
	13'h0860: q2 = 16'h0001; // 0x10c0
	13'h0861: q2 = 16'h81fc; // 0x10c2
	13'h0862: q2 = 16'h9079; // 0x10c4
	13'h0863: q2 = 16'h0001; // 0x10c6
	13'h0864: q2 = 16'h7fb6; // 0x10c8
	13'h0865: q2 = 16'h33c0; // 0x10ca
	13'h0866: q2 = 16'h0001; // 0x10cc
	13'h0867: q2 = 16'h81fc; // 0x10ce
	13'h0868: q2 = 16'h4e5e; // 0x10d0
	13'h0869: q2 = 16'h4e75; // 0x10d2
	13'h086a: q2 = 16'h4e56; // 0x10d4
	13'h086b: q2 = 16'hfffc; // 0x10d6
	13'h086c: q2 = 16'h33fc; // 0x10d8
	13'h086d: q2 = 16'h0001; // 0x10da
	13'h086e: q2 = 16'h0001; // 0x10dc
	13'h086f: q2 = 16'h7fb6; // 0x10de
	13'h0870: q2 = 16'h33fc; // 0x10e0
	13'h0871: q2 = 16'h0020; // 0x10e2
	13'h0872: q2 = 16'h0001; // 0x10e4
	13'h0873: q2 = 16'h81fc; // 0x10e6
	13'h0874: q2 = 16'h4e5e; // 0x10e8
	13'h0875: q2 = 16'h4e75; // 0x10ea
	13'h0876: q2 = 16'h4e56; // 0x10ec
	13'h0877: q2 = 16'hfffc; // 0x10ee
	13'h0878: q2 = 16'h4279; // 0x10f0
	13'h0879: q2 = 16'h0001; // 0x10f2
	13'h087a: q2 = 16'h7fb6; // 0x10f4
	13'h087b: q2 = 16'h4e5e; // 0x10f6
	13'h087c: q2 = 16'h4e75; // 0x10f8
	13'h087d: q2 = 16'h4e56; // 0x10fa
	13'h087e: q2 = 16'hffd2; // 0x10fc
	13'h087f: q2 = 16'h48e7; // 0x10fe
	13'h0880: q2 = 16'h3f1c; // 0x1100
	13'h0881: q2 = 16'h287c; // 0x1102
	13'h0882: q2 = 16'h0001; // 0x1104
	13'h0883: q2 = 16'h75e8; // 0x1106
	13'h0884: q2 = 16'h3e2e; // 0x1108
	13'h0885: q2 = 16'h000a; // 0x110a
	13'h0886: q2 = 16'hde6e; // 0x110c
	13'h0887: q2 = 16'h0008; // 0x110e
	13'h0888: q2 = 16'h5347; // 0x1110
	13'h0889: q2 = 16'h4a79; // 0x1112
	13'h088a: q2 = 16'h0001; // 0x1114
	13'h088b: q2 = 16'h7586; // 0x1116
	13'h088c: q2 = 16'h6700; // 0x1118
	13'h088d: q2 = 16'h008e; // 0x111a
	13'h088e: q2 = 16'h3039; // 0x111c
	13'h088f: q2 = 16'h0001; // 0x111e
	13'h0890: q2 = 16'h7fc0; // 0x1120
	13'h0891: q2 = 16'he340; // 0x1122
	13'h0892: q2 = 16'h48c0; // 0x1124
	13'h0893: q2 = 16'hd0bc; // 0x1126
	13'h0894: q2 = 16'h0000; // 0x1128
	13'h0895: q2 = 16'hf94e; // 0x112a
	13'h0896: q2 = 16'h2040; // 0x112c
	13'h0897: q2 = 16'h3010; // 0x112e
	13'h0898: q2 = 16'hb047; // 0x1130
	13'h0899: q2 = 16'h6e08; // 0x1132
	13'h089a: q2 = 16'h5279; // 0x1134
	13'h089b: q2 = 16'h0001; // 0x1136
	13'h089c: q2 = 16'h7fc0; // 0x1138
	13'h089d: q2 = 16'h601e; // 0x113a
	13'h089e: q2 = 16'h3039; // 0x113c
	13'h089f: q2 = 16'h0001; // 0x113e
	13'h08a0: q2 = 16'h7fc0; // 0x1140
	13'h08a1: q2 = 16'he340; // 0x1142
	13'h08a2: q2 = 16'h48c0; // 0x1144
	13'h08a3: q2 = 16'hd0bc; // 0x1146
	13'h08a4: q2 = 16'h0000; // 0x1148
	13'h08a5: q2 = 16'hf94c; // 0x114a
	13'h08a6: q2 = 16'h2040; // 0x114c
	13'h08a7: q2 = 16'h3010; // 0x114e
	13'h08a8: q2 = 16'hb047; // 0x1150
	13'h08a9: q2 = 16'h6f06; // 0x1152
	13'h08aa: q2 = 16'h5379; // 0x1154
	13'h08ab: q2 = 16'h0001; // 0x1156
	13'h08ac: q2 = 16'h7fc0; // 0x1158
	13'h08ad: q2 = 16'h2079; // 0x115a
	13'h08ae: q2 = 16'h0001; // 0x115c
	13'h08af: q2 = 16'h7fb8; // 0x115e
	13'h08b0: q2 = 16'h3239; // 0x1160
	13'h08b1: q2 = 16'h0001; // 0x1162
	13'h08b2: q2 = 16'h7fce; // 0x1164
	13'h08b3: q2 = 16'hd279; // 0x1166
	13'h08b4: q2 = 16'h0001; // 0x1168
	13'h08b5: q2 = 16'h7fc0; // 0x116a
	13'h08b6: q2 = 16'h5241; // 0x116c
	13'h08b7: q2 = 16'h3141; // 0x116e
	13'h08b8: q2 = 16'h0002; // 0x1170
	13'h08b9: q2 = 16'h3ebc; // 0x1172
	13'h08ba: q2 = 16'h0010; // 0x1174
	13'h08bb: q2 = 16'h4eb9; // 0x1176
	13'h08bc: q2 = 16'h0000; // 0x1178
	13'h08bd: q2 = 16'h549c; // 0x117a
	13'h08be: q2 = 16'h2079; // 0x117c
	13'h08bf: q2 = 16'h0001; // 0x117e
	13'h08c0: q2 = 16'h7fb8; // 0x1180
	13'h08c1: q2 = 16'h5368; // 0x1182
	13'h08c2: q2 = 16'h0002; // 0x1184
	13'h08c3: q2 = 16'h426e; // 0x1186
	13'h08c4: q2 = 16'hffd6; // 0x1188
	13'h08c5: q2 = 16'h302e; // 0x118a
	13'h08c6: q2 = 16'hffd6; // 0x118c
	13'h08c7: q2 = 16'he340; // 0x118e
	13'h08c8: q2 = 16'h48c0; // 0x1190
	13'h08c9: q2 = 16'hd0bc; // 0x1192
	13'h08ca: q2 = 16'h0000; // 0x1194
	13'h08cb: q2 = 16'hf94e; // 0x1196
	13'h08cc: q2 = 16'h2040; // 0x1198
	13'h08cd: q2 = 16'h3010; // 0x119a
	13'h08ce: q2 = 16'hb06e; // 0x119c
	13'h08cf: q2 = 16'h000a; // 0x119e
	13'h08d0: q2 = 16'h6e06; // 0x11a0
	13'h08d1: q2 = 16'h526e; // 0x11a2
	13'h08d2: q2 = 16'hffd6; // 0x11a4
	13'h08d3: q2 = 16'h60e2; // 0x11a6
	13'h08d4: q2 = 16'h4a6e; // 0x11a8
	13'h08d5: q2 = 16'h000c; // 0x11aa
	13'h08d6: q2 = 16'h6f34; // 0x11ac
	13'h08d7: q2 = 16'h4bec; // 0x11ae
	13'h08d8: q2 = 16'h01a2; // 0x11b0
	13'h08d9: q2 = 16'h4246; // 0x11b2
	13'h08da: q2 = 16'hbc7c; // 0x11b4
	13'h08db: q2 = 16'h0009; // 0x11b6
	13'h08dc: q2 = 16'h6c18; // 0x11b8
	13'h08dd: q2 = 16'h7a01; // 0x11ba
	13'h08de: q2 = 16'hba7c; // 0x11bc
	13'h08df: q2 = 16'h0003; // 0x11be
	13'h08e0: q2 = 16'h6e0a; // 0x11c0
	13'h08e1: q2 = 16'h3aad; // 0x11c2
	13'h08e2: q2 = 16'h0008; // 0x11c4
	13'h08e3: q2 = 16'h5245; // 0x11c6
	13'h08e4: q2 = 16'h548d; // 0x11c8
	13'h08e5: q2 = 16'h60f0; // 0x11ca
	13'h08e6: q2 = 16'h548d; // 0x11cc
	13'h08e7: q2 = 16'h5246; // 0x11ce
	13'h08e8: q2 = 16'h60e2; // 0x11d0
	13'h08e9: q2 = 16'h302e; // 0x11d2
	13'h08ea: q2 = 16'h000a; // 0x11d4
	13'h08eb: q2 = 16'hd07c; // 0x11d6
	13'h08ec: q2 = 16'h000a; // 0x11d8
	13'h08ed: q2 = 16'h5340; // 0x11da
	13'h08ee: q2 = 16'h3d40; // 0x11dc
	13'h08ef: q2 = 16'hfffe; // 0x11de
	13'h08f0: q2 = 16'h783d; // 0x11e0
	13'h08f1: q2 = 16'h4a6e; // 0x11e2
	13'h08f2: q2 = 16'h000c; // 0x11e4
	13'h08f3: q2 = 16'h6c2e; // 0x11e6
	13'h08f4: q2 = 16'h4bec; // 0x11e8
	13'h08f5: q2 = 16'h01ee; // 0x11ea
	13'h08f6: q2 = 16'h7c09; // 0x11ec
	13'h08f7: q2 = 16'h4a46; // 0x11ee
	13'h08f8: q2 = 16'h6f1c; // 0x11f0
	13'h08f9: q2 = 16'h7a03; // 0x11f2
	13'h08fa: q2 = 16'hba7c; // 0x11f4
	13'h08fb: q2 = 16'h0001; // 0x11f6
	13'h08fc: q2 = 16'h6d0e; // 0x11f8
	13'h08fd: q2 = 16'h200d; // 0x11fa
	13'h08fe: q2 = 16'h5180; // 0x11fc
	13'h08ff: q2 = 16'h2040; // 0x11fe
	13'h0900: q2 = 16'h3a90; // 0x1200
	13'h0901: q2 = 16'h5345; // 0x1202
	13'h0902: q2 = 16'h558d; // 0x1204
	13'h0903: q2 = 16'h60ec; // 0x1206
	13'h0904: q2 = 16'h558d; // 0x1208
	13'h0905: q2 = 16'h5346; // 0x120a
	13'h0906: q2 = 16'h60e0; // 0x120c
	13'h0907: q2 = 16'h3d6e; // 0x120e
	13'h0908: q2 = 16'h000a; // 0x1210
	13'h0909: q2 = 16'hfffe; // 0x1212
	13'h090a: q2 = 16'h7834; // 0x1214
	13'h090b: q2 = 16'h4a6e; // 0x1216
	13'h090c: q2 = 16'h000c; // 0x1218
	13'h090d: q2 = 16'h6724; // 0x121a
	13'h090e: q2 = 16'h3e84; // 0x121c
	13'h090f: q2 = 16'h200e; // 0x121e
	13'h0910: q2 = 16'hd0bc; // 0x1220
	13'h0911: q2 = 16'hffff; // 0x1222
	13'h0912: q2 = 16'hfff4; // 0x1224
	13'h0913: q2 = 16'h2f00; // 0x1226
	13'h0914: q2 = 16'h200e; // 0x1228
	13'h0915: q2 = 16'hd0bc; // 0x122a
	13'h0916: q2 = 16'hffff; // 0x122c
	13'h0917: q2 = 16'hfffa; // 0x122e
	13'h0918: q2 = 16'h2f00; // 0x1230
	13'h0919: q2 = 16'h3f2e; // 0x1232
	13'h091a: q2 = 16'hfffe; // 0x1234
	13'h091b: q2 = 16'h4eb9; // 0x1236
	13'h091c: q2 = 16'h0000; // 0x1238
	13'h091d: q2 = 16'h1402; // 0x123a
	13'h091e: q2 = 16'hdefc; // 0x123c
	13'h091f: q2 = 16'h000a; // 0x123e
	13'h0920: q2 = 16'h3ebc; // 0x1240
	13'h0921: q2 = 16'h0020; // 0x1242
	13'h0922: q2 = 16'h200e; // 0x1244
	13'h0923: q2 = 16'hd0bc; // 0x1246
	13'h0924: q2 = 16'hffff; // 0x1248
	13'h0925: q2 = 16'hfff4; // 0x124a
	13'h0926: q2 = 16'h2f00; // 0x124c
	13'h0927: q2 = 16'h200e; // 0x124e
	13'h0928: q2 = 16'hd0bc; // 0x1250
	13'h0929: q2 = 16'hffff; // 0x1252
	13'h092a: q2 = 16'hfffa; // 0x1254
	13'h092b: q2 = 16'h2f00; // 0x1256
	13'h092c: q2 = 16'h3f07; // 0x1258
	13'h092d: q2 = 16'h4eb9; // 0x125a
	13'h092e: q2 = 16'h0000; // 0x125c
	13'h092f: q2 = 16'h1402; // 0x125e
	13'h0930: q2 = 16'hdefc; // 0x1260
	13'h0931: q2 = 16'h000a; // 0x1262
	13'h0932: q2 = 16'h302e; // 0x1264
	13'h0933: q2 = 16'hfffa; // 0x1266
	13'h0934: q2 = 16'h5340; // 0x1268
	13'h0935: q2 = 16'he340; // 0x126a
	13'h0936: q2 = 16'h48c0; // 0x126c
	13'h0937: q2 = 16'hd08e; // 0x126e
	13'h0938: q2 = 16'h2040; // 0x1270
	13'h0939: q2 = 16'h3968; // 0x1272
	13'h093a: q2 = 16'hfff4; // 0x1274
	13'h093b: q2 = 16'h010a; // 0x1276
	13'h093c: q2 = 16'h3e87; // 0x1278
	13'h093d: q2 = 16'h4eb9; // 0x127a
	13'h093e: q2 = 16'h0000; // 0x127c
	13'h093f: q2 = 16'h14d0; // 0x127e
	13'h0940: q2 = 16'h4257; // 0x1280
	13'h0941: q2 = 16'h4eb9; // 0x1282
	13'h0942: q2 = 16'h0000; // 0x1284
	13'h0943: q2 = 16'h8a22; // 0x1286
	13'h0944: q2 = 16'h3ebc; // 0x1288
	13'h0945: q2 = 16'h000a; // 0x128a
	13'h0946: q2 = 16'h200e; // 0x128c
	13'h0947: q2 = 16'hd0bc; // 0x128e
	13'h0948: q2 = 16'hffff; // 0x1290
	13'h0949: q2 = 16'hffd8; // 0x1292
	13'h094a: q2 = 16'h2f00; // 0x1294
	13'h094b: q2 = 16'h4eb9; // 0x1296
	13'h094c: q2 = 16'h0000; // 0x1298
	13'h094d: q2 = 16'h78f6; // 0x129a
	13'h094e: q2 = 16'h4a9f; // 0x129c
	13'h094f: q2 = 16'h200e; // 0x129e
	13'h0950: q2 = 16'hd0bc; // 0x12a0
	13'h0951: q2 = 16'hffff; // 0x12a2
	13'h0952: q2 = 16'hffd8; // 0x12a4
	13'h0953: q2 = 16'h2e80; // 0x12a6
	13'h0954: q2 = 16'h4eb9; // 0x12a8
	13'h0955: q2 = 16'h0000; // 0x12aa
	13'h0956: q2 = 16'h072e; // 0x12ac
	13'h0957: q2 = 16'h3a00; // 0x12ae
	13'h0958: q2 = 16'h200e; // 0x12b0
	13'h0959: q2 = 16'hd0bc; // 0x12b2
	13'h095a: q2 = 16'hffff; // 0x12b4
	13'h095b: q2 = 16'hffd8; // 0x12b6
	13'h095c: q2 = 16'h2e80; // 0x12b8
	13'h095d: q2 = 16'h3f07; // 0x12ba
	13'h095e: q2 = 16'h4eb9; // 0x12bc
	13'h095f: q2 = 16'h0000; // 0x12be
	13'h0960: q2 = 16'h0828; // 0x12c0
	13'h0961: q2 = 16'h4a5f; // 0x12c2
	13'h0962: q2 = 16'h7c01; // 0x12c4
	13'h0963: q2 = 16'hbc6e; // 0x12c6
	13'h0964: q2 = 16'hfffa; // 0x12c8
	13'h0965: q2 = 16'h6e32; // 0x12ca
	13'h0966: q2 = 16'h3e86; // 0x12cc
	13'h0967: q2 = 16'h0657; // 0x12ce
	13'h0968: q2 = 16'h0021; // 0x12d0
	13'h0969: q2 = 16'h3006; // 0x12d2
	13'h096a: q2 = 16'h5340; // 0x12d4
	13'h096b: q2 = 16'h48c0; // 0x12d6
	13'h096c: q2 = 16'hd08e; // 0x12d8
	13'h096d: q2 = 16'h2040; // 0x12da
	13'h096e: q2 = 16'h1028; // 0x12dc
	13'h096f: q2 = 16'hffd8; // 0x12de
	13'h0970: q2 = 16'h4880; // 0x12e0
	13'h0971: q2 = 16'h3f00; // 0x12e2
	13'h0972: q2 = 16'h3f3c; // 0x12e4
	13'h0973: q2 = 16'h0012; // 0x12e6
	13'h0974: q2 = 16'h3f05; // 0x12e8
	13'h0975: q2 = 16'h3006; // 0x12ea
	13'h0976: q2 = 16'hd157; // 0x12ec
	13'h0977: q2 = 16'h0657; // 0x12ee
	13'h0978: q2 = 16'h000f; // 0x12f0
	13'h0979: q2 = 16'h4eb9; // 0x12f2
	13'h097a: q2 = 16'h0000; // 0x12f4
	13'h097b: q2 = 16'h3d18; // 0x12f6
	13'h097c: q2 = 16'h5c4f; // 0x12f8
	13'h097d: q2 = 16'h5246; // 0x12fa
	13'h097e: q2 = 16'h60c8; // 0x12fc
	13'h097f: q2 = 16'h7019; // 0x12fe
	13'h0980: q2 = 16'h7203; // 0x1300
	13'h0981: q2 = 16'h926e; // 0x1302
	13'h0982: q2 = 16'hfffa; // 0x1304
	13'h0983: q2 = 16'h9041; // 0x1306
	13'h0984: q2 = 16'h3a00; // 0x1308
	13'h0985: q2 = 16'h7801; // 0x130a
	13'h0986: q2 = 16'h7c19; // 0x130c
	13'h0987: q2 = 16'hbc7c; // 0x130e
	13'h0988: q2 = 16'h0015; // 0x1310
	13'h0989: q2 = 16'h6d64; // 0x1312
	13'h098a: q2 = 16'hbc45; // 0x1314
	13'h098b: q2 = 16'h6634; // 0x1316
	13'h098c: q2 = 16'hb86e; // 0x1318
	13'h098d: q2 = 16'hfffa; // 0x131a
	13'h098e: q2 = 16'h6e2e; // 0x131c
	13'h098f: q2 = 16'h3004; // 0x131e
	13'h0990: q2 = 16'h5340; // 0x1320
	13'h0991: q2 = 16'h48c0; // 0x1322
	13'h0992: q2 = 16'hd08e; // 0x1324
	13'h0993: q2 = 16'h2040; // 0x1326
	13'h0994: q2 = 16'h1028; // 0x1328
	13'h0995: q2 = 16'hffd8; // 0x132a
	13'h0996: q2 = 16'h4880; // 0x132c
	13'h0997: q2 = 16'h3e80; // 0x132e
	13'h0998: q2 = 16'h0657; // 0x1330
	13'h0999: q2 = 16'hffd0; // 0x1332
	13'h099a: q2 = 16'h200e; // 0x1334
	13'h099b: q2 = 16'hd0bc; // 0x1336
	13'h099c: q2 = 16'hffff; // 0x1338
	13'h099d: q2 = 16'hffdc; // 0x133a
	13'h099e: q2 = 16'h2f00; // 0x133c
	13'h099f: q2 = 16'h4eb9; // 0x133e
	13'h09a0: q2 = 16'h0000; // 0x1340
	13'h09a1: q2 = 16'h78f6; // 0x1342
	13'h09a2: q2 = 16'h4a9f; // 0x1344
	13'h09a3: q2 = 16'h5545; // 0x1346
	13'h09a4: q2 = 16'h5244; // 0x1348
	13'h09a5: q2 = 16'h6004; // 0x134a
	13'h09a6: q2 = 16'h422e; // 0x134c
	13'h09a7: q2 = 16'hffdc; // 0x134e
	13'h09a8: q2 = 16'h3e84; // 0x1350
	13'h09a9: q2 = 16'h0657; // 0x1352
	13'h09aa: q2 = 16'h0020; // 0x1354
	13'h09ab: q2 = 16'h3f3c; // 0x1356
	13'h09ac: q2 = 16'h0011; // 0x1358
	13'h09ad: q2 = 16'h3f3c; // 0x135a
	13'h09ae: q2 = 16'h000f; // 0x135c
	13'h09af: q2 = 16'h3f06; // 0x135e
	13'h09b0: q2 = 16'h200e; // 0x1360
	13'h09b1: q2 = 16'hd0bc; // 0x1362
	13'h09b2: q2 = 16'hffff; // 0x1364
	13'h09b3: q2 = 16'hffdc; // 0x1366
	13'h09b4: q2 = 16'h2f00; // 0x1368
	13'h09b5: q2 = 16'h4eb9; // 0x136a
	13'h09b6: q2 = 16'h0000; // 0x136c
	13'h09b7: q2 = 16'h026c; // 0x136e
	13'h09b8: q2 = 16'hdefc; // 0x1370
	13'h09b9: q2 = 16'h000a; // 0x1372
	13'h09ba: q2 = 16'h5346; // 0x1374
	13'h09bb: q2 = 16'h6096; // 0x1376
	13'h09bc: q2 = 16'hbe7c; // 0x1378
	13'h09bd: q2 = 16'h000a; // 0x137a
	13'h09be: q2 = 16'h6c08; // 0x137c
	13'h09bf: q2 = 16'h267c; // 0x137e
	13'h09c0: q2 = 16'h0000; // 0x1380
	13'h09c1: q2 = 16'hc556; // 0x1382
	13'h09c2: q2 = 16'h6014; // 0x1384
	13'h09c3: q2 = 16'hbe7c; // 0x1386
	13'h09c4: q2 = 16'h0064; // 0x1388
	13'h09c5: q2 = 16'h6c08; // 0x138a
	13'h09c6: q2 = 16'h267c; // 0x138c
	13'h09c7: q2 = 16'h0000; // 0x138e
	13'h09c8: q2 = 16'hc59e; // 0x1390
	13'h09c9: q2 = 16'h6006; // 0x1392
	13'h09ca: q2 = 16'h267c; // 0x1394
	13'h09cb: q2 = 16'h0000; // 0x1396
	13'h09cc: q2 = 16'hc5e6; // 0x1398
	13'h09cd: q2 = 16'h7c03; // 0x139a
	13'h09ce: q2 = 16'hbc7c; // 0x139c
	13'h09cf: q2 = 16'h000c; // 0x139e
	13'h09d0: q2 = 16'h6c40; // 0x13a0
	13'h09d1: q2 = 16'h7a1a; // 0x13a2
	13'h09d2: q2 = 16'hba7c; // 0x13a4
	13'h09d3: q2 = 16'h0013; // 0x13a6
	13'h09d4: q2 = 16'h6d34; // 0x13a8
	13'h09d5: q2 = 16'h1013; // 0x13aa
	13'h09d6: q2 = 16'h4880; // 0x13ac
	13'h09d7: q2 = 16'hc07c; // 0x13ae
	13'h09d8: q2 = 16'h00ff; // 0x13b0
	13'h09d9: q2 = 16'h3d40; // 0x13b2
	13'h09da: q2 = 16'hfffc; // 0x13b4
	13'h09db: q2 = 16'h0c6e; // 0x13b6
	13'h09dc: q2 = 16'h0020; // 0x13b8
	13'h09dd: q2 = 16'hfffc; // 0x13ba
	13'h09de: q2 = 16'h6c06; // 0x13bc
	13'h09df: q2 = 16'h066e; // 0x13be
	13'h09e0: q2 = 16'h0100; // 0x13c0
	13'h09e1: q2 = 16'hfffc; // 0x13c2
	13'h09e2: q2 = 16'h3ebc; // 0x13c4
	13'h09e3: q2 = 16'h0020; // 0x13c6
	13'h09e4: q2 = 16'h3f2e; // 0x13c8
	13'h09e5: q2 = 16'hfffc; // 0x13ca
	13'h09e6: q2 = 16'h3f05; // 0x13cc
	13'h09e7: q2 = 16'h3f06; // 0x13ce
	13'h09e8: q2 = 16'h4eb9; // 0x13d0
	13'h09e9: q2 = 16'h0000; // 0x13d2
	13'h09ea: q2 = 16'h3d18; // 0x13d4
	13'h09eb: q2 = 16'h5c4f; // 0x13d6
	13'h09ec: q2 = 16'h528b; // 0x13d8
	13'h09ed: q2 = 16'h5345; // 0x13da
	13'h09ee: q2 = 16'h60c6; // 0x13dc
	13'h09ef: q2 = 16'h5246; // 0x13de
	13'h09f0: q2 = 16'h60ba; // 0x13e0
	13'h09f1: q2 = 16'h7834; // 0x13e2
	13'h09f2: q2 = 16'h3d6e; // 0x13e4
	13'h09f3: q2 = 16'h000a; // 0x13e6
	13'h09f4: q2 = 16'hfffe; // 0x13e8
	13'h09f5: q2 = 16'h3d6e; // 0x13ea
	13'h09f6: q2 = 16'hffd6; // 0x13ec
	13'h09f7: q2 = 16'hffd4; // 0x13ee
	13'h09f8: q2 = 16'h3d7c; // 0x13f0
	13'h09f9: q2 = 16'h0002; // 0x13f2
	13'h09fa: q2 = 16'hffee; // 0x13f4
	13'h09fb: q2 = 16'h362e; // 0x13f6
	13'h09fc: q2 = 16'hffee; // 0x13f8
	13'h09fd: q2 = 16'h4246; // 0x13fa
	13'h09fe: q2 = 16'hbc7c; // 0x13fc
	13'h09ff: q2 = 16'h000a; // 0x13fe
	13'h0a00: q2 = 16'h6c00; // 0x1400
	13'h0a01: q2 = 16'h0164; // 0x1402
	13'h0a02: q2 = 16'h0c6e; // 0x1404
	13'h0a03: q2 = 16'h000a; // 0x1406
	13'h0a04: q2 = 16'hfffe; // 0x1408
	13'h0a05: q2 = 16'h6c08; // 0x140a
	13'h0a06: q2 = 16'h3d7c; // 0x140c
	13'h0a07: q2 = 16'h00e9; // 0x140e
	13'h0a08: q2 = 16'hfffc; // 0x1410
	13'h0a09: q2 = 16'h6016; // 0x1412
	13'h0a0a: q2 = 16'h0c6e; // 0x1414
	13'h0a0b: q2 = 16'h0064; // 0x1416
	13'h0a0c: q2 = 16'hfffe; // 0x1418
	13'h0a0d: q2 = 16'h6c08; // 0x141a
	13'h0a0e: q2 = 16'h3d7c; // 0x141c
	13'h0a0f: q2 = 16'h00e1; // 0x141e
	13'h0a10: q2 = 16'hfffc; // 0x1420
	13'h0a11: q2 = 16'h6006; // 0x1422
	13'h0a12: q2 = 16'h3d7c; // 0x1424
	13'h0a13: q2 = 16'h00d9; // 0x1426
	13'h0a14: q2 = 16'hfffc; // 0x1428
	13'h0a15: q2 = 16'h3e84; // 0x142a
	13'h0a16: q2 = 16'h3f2e; // 0x142c
	13'h0a17: q2 = 16'hfffc; // 0x142e
	13'h0a18: q2 = 16'h3f3c; // 0x1430
	13'h0a19: q2 = 16'h000a; // 0x1432
	13'h0a1a: q2 = 16'h3f03; // 0x1434
	13'h0a1b: q2 = 16'h4eb9; // 0x1436
	13'h0a1c: q2 = 16'h0000; // 0x1438
	13'h0a1d: q2 = 16'h3d18; // 0x143a
	13'h0a1e: q2 = 16'h5c4f; // 0x143c
	13'h0a1f: q2 = 16'h302e; // 0x143e
	13'h0a20: q2 = 16'hfffe; // 0x1440
	13'h0a21: q2 = 16'h48c0; // 0x1442
	13'h0a22: q2 = 16'h81fc; // 0x1444
	13'h0a23: q2 = 16'h0005; // 0x1446
	13'h0a24: q2 = 16'h4840; // 0x1448
	13'h0a25: q2 = 16'h4a40; // 0x144a
	13'h0a26: q2 = 16'h6610; // 0x144c
	13'h0a27: q2 = 16'h0c6e; // 0x144e
	13'h0a28: q2 = 16'h007d; // 0x1450
	13'h0a29: q2 = 16'hfffe; // 0x1452
	13'h0a2a: q2 = 16'h6708; // 0x1454
	13'h0a2b: q2 = 16'h3d7c; // 0x1456
	13'h0a2c: q2 = 16'h0018; // 0x1458
	13'h0a2d: q2 = 16'hffd2; // 0x145a
	13'h0a2e: q2 = 16'h6004; // 0x145c
	13'h0a2f: q2 = 16'h426e; // 0x145e
	13'h0a30: q2 = 16'hffd2; // 0x1460
	13'h0a31: q2 = 16'h3d7c; // 0x1462
	13'h0a32: q2 = 16'h0008; // 0x1464
	13'h0a33: q2 = 16'hfff0; // 0x1466
	13'h0a34: q2 = 16'h3003; // 0x1468
	13'h0a35: q2 = 16'h5340; // 0x146a
	13'h0a36: q2 = 16'h3d40; // 0x146c
	13'h0a37: q2 = 16'hfff2; // 0x146e
	13'h0a38: q2 = 16'h7a66; // 0x1470
	13'h0a39: q2 = 16'hba7c; // 0x1472
	13'h0a3a: q2 = 16'h006b; // 0x1474
	13'h0a3b: q2 = 16'h6e34; // 0x1476
	13'h0a3c: q2 = 16'h3eae; // 0x1478
	13'h0a3d: q2 = 16'hffd2; // 0x147a
	13'h0a3e: q2 = 16'h3f05; // 0x147c
	13'h0a3f: q2 = 16'h3f2e; // 0x147e
	13'h0a40: q2 = 16'hfff0; // 0x1480
	13'h0a41: q2 = 16'h3f2e; // 0x1482
	13'h0a42: q2 = 16'hfff2; // 0x1484
	13'h0a43: q2 = 16'h4eb9; // 0x1486
	13'h0a44: q2 = 16'h0000; // 0x1488
	13'h0a45: q2 = 16'h3d18; // 0x148a
	13'h0a46: q2 = 16'h5c4f; // 0x148c
	13'h0a47: q2 = 16'h526e; // 0x148e
	13'h0a48: q2 = 16'hfff2; // 0x1490
	13'h0a49: q2 = 16'h3003; // 0x1492
	13'h0a4a: q2 = 16'h5240; // 0x1494
	13'h0a4b: q2 = 16'hb06e; // 0x1496
	13'h0a4c: q2 = 16'hfff2; // 0x1498
	13'h0a4d: q2 = 16'h6c0c; // 0x149a
	13'h0a4e: q2 = 16'h3003; // 0x149c
	13'h0a4f: q2 = 16'h5340; // 0x149e
	13'h0a50: q2 = 16'h3d40; // 0x14a0
	13'h0a51: q2 = 16'hfff2; // 0x14a2
	13'h0a52: q2 = 16'h536e; // 0x14a4
	13'h0a53: q2 = 16'hfff0; // 0x14a6
	13'h0a54: q2 = 16'h5245; // 0x14a8
	13'h0a55: q2 = 16'h60c6; // 0x14aa
	13'h0a56: q2 = 16'h0c6e; // 0x14ac
	13'h0a57: q2 = 16'h007d; // 0x14ae
	13'h0a58: q2 = 16'hfffe; // 0x14b0
	13'h0a59: q2 = 16'h6616; // 0x14b2
	13'h0a5a: q2 = 16'h3ebc; // 0x14b4
	13'h0a5b: q2 = 16'h003e; // 0x14b6
	13'h0a5c: q2 = 16'h3f3c; // 0x14b8
	13'h0a5d: q2 = 16'h003f; // 0x14ba
	13'h0a5e: q2 = 16'h3f3c; // 0x14bc
	13'h0a5f: q2 = 16'h0007; // 0x14be
	13'h0a60: q2 = 16'h3f03; // 0x14c0
	13'h0a61: q2 = 16'h4eb9; // 0x14c2
	13'h0a62: q2 = 16'h0000; // 0x14c4
	13'h0a63: q2 = 16'h3d18; // 0x14c6
	13'h0a64: q2 = 16'h5c4f; // 0x14c8
	13'h0a65: q2 = 16'h4a79; // 0x14ca
	13'h0a66: q2 = 16'h0001; // 0x14cc
	13'h0a67: q2 = 16'h7586; // 0x14ce
	13'h0a68: q2 = 16'h6724; // 0x14d0
	13'h0a69: q2 = 16'h302e; // 0x14d2
	13'h0a6a: q2 = 16'hffd4; // 0x14d4
	13'h0a6b: q2 = 16'he340; // 0x14d6
	13'h0a6c: q2 = 16'h48c0; // 0x14d8
	13'h0a6d: q2 = 16'hd0bc; // 0x14da
	13'h0a6e: q2 = 16'h0000; // 0x14dc
	13'h0a6f: q2 = 16'hf94e; // 0x14de
	13'h0a70: q2 = 16'h2040; // 0x14e0
	13'h0a71: q2 = 16'h3010; // 0x14e2
	13'h0a72: q2 = 16'hb06e; // 0x14e4
	13'h0a73: q2 = 16'hfffe; // 0x14e6
	13'h0a74: q2 = 16'h6e0c; // 0x14e8
	13'h0a75: q2 = 16'h526e; // 0x14ea
	13'h0a76: q2 = 16'hffd4; // 0x14ec
	13'h0a77: q2 = 16'h3d7c; // 0x14ee
	13'h0a78: q2 = 16'h0007; // 0x14f0
	13'h0a79: q2 = 16'hfff0; // 0x14f2
	13'h0a7a: q2 = 16'h6004; // 0x14f4
	13'h0a7b: q2 = 16'h426e; // 0x14f6
	13'h0a7c: q2 = 16'hfff0; // 0x14f8
	13'h0a7d: q2 = 16'h426e; // 0x14fa
	13'h0a7e: q2 = 16'hfff2; // 0x14fc
	13'h0a7f: q2 = 16'h7a14; // 0x14fe
	13'h0a80: q2 = 16'hba7c; // 0x1500
	13'h0a81: q2 = 16'h0015; // 0x1502
	13'h0a82: q2 = 16'h6e30; // 0x1504
	13'h0a83: q2 = 16'h3eae; // 0x1506
	13'h0a84: q2 = 16'hfff0; // 0x1508
	13'h0a85: q2 = 16'h3f05; // 0x150a
	13'h0a86: q2 = 16'h3f3c; // 0x150c
	13'h0a87: q2 = 16'h0006; // 0x150e
	13'h0a88: q2 = 16'h3f03; // 0x1510
	13'h0a89: q2 = 16'h302e; // 0x1512
	13'h0a8a: q2 = 16'hfff2; // 0x1514
	13'h0a8b: q2 = 16'hd157; // 0x1516
	13'h0a8c: q2 = 16'h4eb9; // 0x1518
	13'h0a8d: q2 = 16'h0000; // 0x151a
	13'h0a8e: q2 = 16'h3d18; // 0x151c
	13'h0a8f: q2 = 16'h5c4f; // 0x151e
	13'h0a90: q2 = 16'h526e; // 0x1520
	13'h0a91: q2 = 16'hfff2; // 0x1522
	13'h0a92: q2 = 16'h0c6e; // 0x1524
	13'h0a93: q2 = 16'h0007; // 0x1526
	13'h0a94: q2 = 16'hfff0; // 0x1528
	13'h0a95: q2 = 16'h6606; // 0x152a
	13'h0a96: q2 = 16'h3d7c; // 0x152c
	13'h0a97: q2 = 16'h002b; // 0x152e
	13'h0a98: q2 = 16'hfff0; // 0x1530
	13'h0a99: q2 = 16'h5245; // 0x1532
	13'h0a9a: q2 = 16'h60ca; // 0x1534
	13'h0a9b: q2 = 16'h302e; // 0x1536
	13'h0a9c: q2 = 16'hfffe; // 0x1538
	13'h0a9d: q2 = 16'hb047; // 0x153a
	13'h0a9e: q2 = 16'h6704; // 0x153c
	13'h0a9f: q2 = 16'h4245; // 0x153e
	13'h0aa0: q2 = 16'h6002; // 0x1540
	13'h0aa1: q2 = 16'h7a3e; // 0x1542
	13'h0aa2: q2 = 16'h3e85; // 0x1544
	13'h0aa3: q2 = 16'h3f3c; // 0x1546
	13'h0aa4: q2 = 16'h006c; // 0x1548
	13'h0aa5: q2 = 16'h3f3c; // 0x154a
	13'h0aa6: q2 = 16'h000b; // 0x154c
	13'h0aa7: q2 = 16'h3f03; // 0x154e
	13'h0aa8: q2 = 16'h4eb9; // 0x1550
	13'h0aa9: q2 = 16'h0000; // 0x1552
	13'h0aaa: q2 = 16'h3d18; // 0x1554
	13'h0aab: q2 = 16'h5c4f; // 0x1556
	13'h0aac: q2 = 16'h5643; // 0x1558
	13'h0aad: q2 = 16'h5244; // 0x155a
	13'h0aae: q2 = 16'h526e; // 0x155c
	13'h0aaf: q2 = 16'hfffe; // 0x155e
	13'h0ab0: q2 = 16'h5246; // 0x1560
	13'h0ab1: q2 = 16'h6000; // 0x1562
	13'h0ab2: q2 = 16'hfe98; // 0x1564
	13'h0ab3: q2 = 16'h4a9f; // 0x1566
	13'h0ab4: q2 = 16'h4cdf; // 0x1568
	13'h0ab5: q2 = 16'h38f8; // 0x156a
	13'h0ab6: q2 = 16'h4e5e; // 0x156c
	13'h0ab7: q2 = 16'h4e75; // 0x156e
	13'h0ab8: q2 = 16'h4e56; // 0x1570
	13'h0ab9: q2 = 16'hffd4; // 0x1572
	13'h0aba: q2 = 16'h48e7; // 0x1574
	13'h0abb: q2 = 16'h3f00; // 0x1576
	13'h0abc: q2 = 16'h4a79; // 0x1578
	13'h0abd: q2 = 16'h0001; // 0x157a
	13'h0abe: q2 = 16'h7588; // 0x157c
	13'h0abf: q2 = 16'h660e; // 0x157e
	13'h0ac0: q2 = 16'h2079; // 0x1580
	13'h0ac1: q2 = 16'h0001; // 0x1582
	13'h0ac2: q2 = 16'h7fb8; // 0x1584
	13'h0ac3: q2 = 16'h4a68; // 0x1586
	13'h0ac4: q2 = 16'h001c; // 0x1588
	13'h0ac5: q2 = 16'h6700; // 0x158a
	13'h0ac6: q2 = 16'h037c; // 0x158c
	13'h0ac7: q2 = 16'h0c79; // 0x158e
	13'h0ac8: q2 = 16'h0003; // 0x1590
	13'h0ac9: q2 = 16'h0001; // 0x1592
	13'h0aca: q2 = 16'h7588; // 0x1594
	13'h0acb: q2 = 16'h660e; // 0x1596
	13'h0acc: q2 = 16'h2079; // 0x1598
	13'h0acd: q2 = 16'h0001; // 0x159a
	13'h0ace: q2 = 16'h7fb8; // 0x159c
	13'h0acf: q2 = 16'h30bc; // 0x159e
	13'h0ad0: q2 = 16'h0001; // 0x15a0
	13'h0ad1: q2 = 16'h6000; // 0x15a2
	13'h0ad2: q2 = 16'h0364; // 0x15a4
	13'h0ad3: q2 = 16'h2a39; // 0x15a6
	13'h0ad4: q2 = 16'h0000; // 0x15a8
	13'h0ad5: q2 = 16'hf96a; // 0x15aa
	13'h0ad6: q2 = 16'h4244; // 0x15ac
	13'h0ad7: q2 = 16'h4eb9; // 0x15ae
	13'h0ad8: q2 = 16'h0000; // 0x15b0
	13'h0ad9: q2 = 16'h0226; // 0x15b2
	13'h0ada: q2 = 16'h2079; // 0x15b4
	13'h0adb: q2 = 16'h0001; // 0x15b6
	13'h0adc: q2 = 16'h7fb8; // 0x15b8
	13'h0add: q2 = 16'h3d50; // 0x15ba
	13'h0ade: q2 = 16'hfff6; // 0x15bc
	13'h0adf: q2 = 16'h0c79; // 0x15be
	13'h0ae0: q2 = 16'h0001; // 0x15c0
	13'h0ae1: q2 = 16'h0001; // 0x15c2
	13'h0ae2: q2 = 16'h7588; // 0x15c4
	13'h0ae3: q2 = 16'h660e; // 0x15c6
	13'h0ae4: q2 = 16'h0c6e; // 0x15c8
	13'h0ae5: q2 = 16'h0009; // 0x15ca
	13'h0ae6: q2 = 16'hfff6; // 0x15cc
	13'h0ae7: q2 = 16'h6c06; // 0x15ce
	13'h0ae8: q2 = 16'h3d7c; // 0x15d0
	13'h0ae9: q2 = 16'h0009; // 0x15d2
	13'h0aea: q2 = 16'hfff6; // 0x15d4
	13'h0aeb: q2 = 16'h0c79; // 0x15d6
	13'h0aec: q2 = 16'h0002; // 0x15d8
	13'h0aed: q2 = 16'h0001; // 0x15da
	13'h0aee: q2 = 16'h7588; // 0x15dc
	13'h0aef: q2 = 16'h6606; // 0x15de
	13'h0af0: q2 = 16'h3d7c; // 0x15e0
	13'h0af1: q2 = 16'h007d; // 0x15e2
	13'h0af2: q2 = 16'hfff6; // 0x15e4
	13'h0af3: q2 = 16'h3d7c; // 0x15e6
	13'h0af4: q2 = 16'h0001; // 0x15e8
	13'h0af5: q2 = 16'hfff8; // 0x15ea
	13'h0af6: q2 = 16'h302e; // 0x15ec
	13'h0af7: q2 = 16'hfff6; // 0x15ee
	13'h0af8: q2 = 16'h5640; // 0x15f0
	13'h0af9: q2 = 16'h3d40; // 0x15f2
	13'h0afa: q2 = 16'hfffa; // 0x15f4
	13'h0afb: q2 = 16'h0c6e; // 0x15f6
	13'h0afc: q2 = 16'h007d; // 0x15f8
	13'h0afd: q2 = 16'hfffa; // 0x15fa
	13'h0afe: q2 = 16'h6f06; // 0x15fc
	13'h0aff: q2 = 16'h3d7c; // 0x15fe
	13'h0b00: q2 = 16'h007d; // 0x1600
	13'h0b01: q2 = 16'hfffa; // 0x1602
	13'h0b02: q2 = 16'h7c01; // 0x1604
	13'h0b03: q2 = 16'h3d7c; // 0x1606
	13'h0b04: q2 = 16'h0001; // 0x1608
	13'h0b05: q2 = 16'hfff4; // 0x160a
	13'h0b06: q2 = 16'h7e01; // 0x160c
	13'h0b07: q2 = 16'h3d7c; // 0x160e
	13'h0b08: q2 = 16'h0001; // 0x1610
	13'h0b09: q2 = 16'hfffe; // 0x1612
	13'h0b0a: q2 = 16'h3d7c; // 0x1614
	13'h0b0b: q2 = 16'h000a; // 0x1616
	13'h0b0c: q2 = 16'hfffc; // 0x1618
	13'h0b0d: q2 = 16'h3d7c; // 0x161a
	13'h0b0e: q2 = 16'h0001; // 0x161c
	13'h0b0f: q2 = 16'hfff2; // 0x161e
	13'h0b10: q2 = 16'h4eb9; // 0x1620
	13'h0b11: q2 = 16'h0000; // 0x1622
	13'h0b12: q2 = 16'h9912; // 0x1624
	13'h0b13: q2 = 16'h4257; // 0x1626
	13'h0b14: q2 = 16'h3f2e; // 0x1628
	13'h0b15: q2 = 16'hfffe; // 0x162a
	13'h0b16: q2 = 16'h3f07; // 0x162c
	13'h0b17: q2 = 16'h4eb9; // 0x162e
	13'h0b18: q2 = 16'h0000; // 0x1630
	13'h0b19: q2 = 16'h90fa; // 0x1632
	13'h0b1a: q2 = 16'h4a9f; // 0x1634
	13'h0b1b: q2 = 16'h23fc; // 0x1636
	13'h0b1c: q2 = 16'h0000; // 0x1638
	13'h0b1d: q2 = 16'h003c; // 0x163a
	13'h0b1e: q2 = 16'h0001; // 0x163c
	13'h0b1f: q2 = 16'h7fc2; // 0x163e
	13'h0b20: q2 = 16'h3d7c; // 0x1640
	13'h0b21: q2 = 16'h000f; // 0x1642
	13'h0b22: q2 = 16'hfff0; // 0x1644
	13'h0b23: q2 = 16'h4a6e; // 0x1646
	13'h0b24: q2 = 16'hfff0; // 0x1648
	13'h0b25: q2 = 16'h6f00; // 0x164a
	13'h0b26: q2 = 16'h0262; // 0x164c
	13'h0b27: q2 = 16'h4ab9; // 0x164e
	13'h0b28: q2 = 16'h0001; // 0x1650
	13'h0b29: q2 = 16'h7fc2; // 0x1652
	13'h0b2a: q2 = 16'h660e; // 0x1654
	13'h0b2b: q2 = 16'h536e; // 0x1656
	13'h0b2c: q2 = 16'hfff0; // 0x1658
	13'h0b2d: q2 = 16'h23fc; // 0x165a
	13'h0b2e: q2 = 16'h0000; // 0x165c
	13'h0b2f: q2 = 16'h003c; // 0x165e
	13'h0b30: q2 = 16'h0001; // 0x1660
	13'h0b31: q2 = 16'h7fc2; // 0x1662
	13'h0b32: q2 = 16'h3ebc; // 0x1664
	13'h0b33: q2 = 16'h000e; // 0x1666
	13'h0b34: q2 = 16'h200e; // 0x1668
	13'h0b35: q2 = 16'hd0bc; // 0x166a
	13'h0b36: q2 = 16'hffff; // 0x166c
	13'h0b37: q2 = 16'hffe4; // 0x166e
	13'h0b38: q2 = 16'h2f00; // 0x1670
	13'h0b39: q2 = 16'h4eb9; // 0x1672
	13'h0b3a: q2 = 16'h0000; // 0x1674
	13'h0b3b: q2 = 16'h78f6; // 0x1676
	13'h0b3c: q2 = 16'h4a9f; // 0x1678
	13'h0b3d: q2 = 16'h0c6e; // 0x167a
	13'h0b3e: q2 = 16'h000a; // 0x167c
	13'h0b3f: q2 = 16'hfff0; // 0x167e
	13'h0b40: q2 = 16'h6c18; // 0x1680
	13'h0b41: q2 = 16'h2ebc; // 0x1682
	13'h0b42: q2 = 16'h0000; // 0x1684
	13'h0b43: q2 = 16'hf97a; // 0x1686
	13'h0b44: q2 = 16'h200e; // 0x1688
	13'h0b45: q2 = 16'hd0bc; // 0x168a
	13'h0b46: q2 = 16'hffff; // 0x168c
	13'h0b47: q2 = 16'hffe4; // 0x168e
	13'h0b48: q2 = 16'h2f00; // 0x1690
	13'h0b49: q2 = 16'h4eb9; // 0x1692
	13'h0b4a: q2 = 16'h0000; // 0x1694
	13'h0b4b: q2 = 16'h0770; // 0x1696
	13'h0b4c: q2 = 16'h4a9f; // 0x1698
	13'h0b4d: q2 = 16'h200e; // 0x169a
	13'h0b4e: q2 = 16'hd0bc; // 0x169c
	13'h0b4f: q2 = 16'hffff; // 0x169e
	13'h0b50: q2 = 16'hffe4; // 0x16a0
	13'h0b51: q2 = 16'h2e80; // 0x16a2
	13'h0b52: q2 = 16'h3f2e; // 0x16a4
	13'h0b53: q2 = 16'hfff0; // 0x16a6
	13'h0b54: q2 = 16'h4eb9; // 0x16a8
	13'h0b55: q2 = 16'h0000; // 0x16aa
	13'h0b56: q2 = 16'h0798; // 0x16ac
	13'h0b57: q2 = 16'h4a5f; // 0x16ae
	13'h0b58: q2 = 16'h3ebc; // 0x16b0
	13'h0b59: q2 = 16'h0031; // 0x16b2
	13'h0b5a: q2 = 16'h3f3c; // 0x16b4
	13'h0b5b: q2 = 16'h000b; // 0x16b6
	13'h0b5c: q2 = 16'h3f3c; // 0x16b8
	13'h0b5d: q2 = 16'hffe3; // 0x16ba
	13'h0b5e: q2 = 16'h3f3c; // 0x16bc
	13'h0b5f: q2 = 16'h000e; // 0x16be
	13'h0b60: q2 = 16'h200e; // 0x16c0
	13'h0b61: q2 = 16'hd0bc; // 0x16c2
	13'h0b62: q2 = 16'hffff; // 0x16c4
	13'h0b63: q2 = 16'hffe4; // 0x16c6
	13'h0b64: q2 = 16'h2f00; // 0x16c8
	13'h0b65: q2 = 16'h4eb9; // 0x16ca
	13'h0b66: q2 = 16'h0000; // 0x16cc
	13'h0b67: q2 = 16'h026c; // 0x16ce
	13'h0b68: q2 = 16'hdefc; // 0x16d0
	13'h0b69: q2 = 16'h000a; // 0x16d2
	13'h0b6a: q2 = 16'h4243; // 0x16d4
	13'h0b6b: q2 = 16'h302e; // 0x16d6
	13'h0b6c: q2 = 16'hfffe; // 0x16d8
	13'h0b6d: q2 = 16'hb06e; // 0x16da
	13'h0b6e: q2 = 16'hfff2; // 0x16dc
	13'h0b6f: q2 = 16'h6f02; // 0x16de
	13'h0b70: q2 = 16'h7601; // 0x16e0
	13'h0b71: q2 = 16'h302e; // 0x16e2
	13'h0b72: q2 = 16'hfffe; // 0x16e4
	13'h0b73: q2 = 16'hb06e; // 0x16e6
	13'h0b74: q2 = 16'hfff2; // 0x16e8
	13'h0b75: q2 = 16'h6c02; // 0x16ea
	13'h0b76: q2 = 16'h76ff; // 0x16ec
	13'h0b77: q2 = 16'hbc6e; // 0x16ee
	13'h0b78: q2 = 16'hfff4; // 0x16f0
	13'h0b79: q2 = 16'h670c; // 0x16f2
	13'h0b7a: q2 = 16'h2ebc; // 0x16f4
	13'h0b7b: q2 = 16'h0000; // 0x16f6
	13'h0b7c: q2 = 16'hfd1c; // 0x16f8
	13'h0b7d: q2 = 16'h4eb9; // 0x16fa
	13'h0b7e: q2 = 16'h0000; // 0x16fc
	13'h0b7f: q2 = 16'h7dd8; // 0x16fe
	13'h0b80: q2 = 16'h3e83; // 0x1700
	13'h0b81: q2 = 16'h3f2e; // 0x1702
	13'h0b82: q2 = 16'hfffe; // 0x1704
	13'h0b83: q2 = 16'h3f07; // 0x1706
	13'h0b84: q2 = 16'h4eb9; // 0x1708
	13'h0b85: q2 = 16'h0000; // 0x170a
	13'h0b86: q2 = 16'h90fa; // 0x170c
	13'h0b87: q2 = 16'h4a9f; // 0x170e
	13'h0b88: q2 = 16'h4a85; // 0x1710
	13'h0b89: q2 = 16'h6f18; // 0x1712
	13'h0b8a: q2 = 16'h23c5; // 0x1714
	13'h0b8b: q2 = 16'h0001; // 0x1716
	13'h0b8c: q2 = 16'h7f60; // 0x1718
	13'h0b8d: q2 = 16'h4ab9; // 0x171a
	13'h0b8e: q2 = 16'h0001; // 0x171c
	13'h0b8f: q2 = 16'h7f60; // 0x171e
	13'h0b90: q2 = 16'h670a; // 0x1720
	13'h0b91: q2 = 16'h4a79; // 0x1722
	13'h0b92: q2 = 16'h0001; // 0x1724
	13'h0b93: q2 = 16'h7fca; // 0x1726
	13'h0b94: q2 = 16'h6602; // 0x1728
	13'h0b95: q2 = 16'h60ee; // 0x172a
	13'h0b96: q2 = 16'h4a79; // 0x172c
	13'h0b97: q2 = 16'h0001; // 0x172e
	13'h0b98: q2 = 16'h7fca; // 0x1730
	13'h0b99: q2 = 16'h6600; // 0x1732
	13'h0b9a: q2 = 16'h017a; // 0x1734
	13'h0b9b: q2 = 16'h3d46; // 0x1736
	13'h0b9c: q2 = 16'hfff4; // 0x1738
	13'h0b9d: q2 = 16'h3d6e; // 0x173a
	13'h0b9e: q2 = 16'hfffe; // 0x173c
	13'h0b9f: q2 = 16'hfff2; // 0x173e
	13'h0ba0: q2 = 16'h302e; // 0x1740
	13'h0ba1: q2 = 16'hfff6; // 0x1742
	13'h0ba2: q2 = 16'h906e; // 0x1744
	13'h0ba3: q2 = 16'hfffe; // 0x1746
	13'h0ba4: q2 = 16'h5240; // 0x1748
	13'h0ba5: q2 = 16'h3d40; // 0x174a
	13'h0ba6: q2 = 16'hffe2; // 0x174c
	13'h0ba7: q2 = 16'h0c6e; // 0x174e
	13'h0ba8: q2 = 16'h007d; // 0x1750
	13'h0ba9: q2 = 16'hfffc; // 0x1752
	13'h0baa: q2 = 16'h670e; // 0x1754
	13'h0bab: q2 = 16'h0c6e; // 0x1756
	13'h0bac: q2 = 16'h0007; // 0x1758
	13'h0bad: q2 = 16'hfff6; // 0x175a
	13'h0bae: q2 = 16'h6d06; // 0x175c
	13'h0baf: q2 = 16'h3d7c; // 0x175e
	13'h0bb0: q2 = 16'h0007; // 0x1760
	13'h0bb1: q2 = 16'hffe2; // 0x1762
	13'h0bb2: q2 = 16'h2079; // 0x1764
	13'h0bb3: q2 = 16'h0001; // 0x1766
	13'h0bb4: q2 = 16'h7eb2; // 0x1768
	13'h0bb5: q2 = 16'h3028; // 0x176a
	13'h0bb6: q2 = 16'h0002; // 0x176c
	13'h0bb7: q2 = 16'h2279; // 0x176e
	13'h0bb8: q2 = 16'h0001; // 0x1770
	13'h0bb9: q2 = 16'h7eb2; // 0x1772
	13'h0bba: q2 = 16'h9051; // 0x1774
	13'h0bbb: q2 = 16'he440; // 0x1776
	13'h0bbc: q2 = 16'h3d40; // 0x1778
	13'h0bbd: q2 = 16'hffe0; // 0x177a
	13'h0bbe: q2 = 16'h302e; // 0x177c
	13'h0bbf: q2 = 16'hffe0; // 0x177e
	13'h0bc0: q2 = 16'h4440; // 0x1780
	13'h0bc1: q2 = 16'hb079; // 0x1782
	13'h0bc2: q2 = 16'h0001; // 0x1784
	13'h0bc3: q2 = 16'h8622; // 0x1786
	13'h0bc4: q2 = 16'h6f08; // 0x1788
	13'h0bc5: q2 = 16'h3d7c; // 0x178a
	13'h0bc6: q2 = 16'h0001; // 0x178c
	13'h0bc7: q2 = 16'hffdc; // 0x178e
	13'h0bc8: q2 = 16'h6004; // 0x1790
	13'h0bc9: q2 = 16'h426e; // 0x1792
	13'h0bca: q2 = 16'hffdc; // 0x1794
	13'h0bcb: q2 = 16'h3039; // 0x1796
	13'h0bcc: q2 = 16'h0001; // 0x1798
	13'h0bcd: q2 = 16'h8622; // 0x179a
	13'h0bce: q2 = 16'hb06e; // 0x179c
	13'h0bcf: q2 = 16'hffe0; // 0x179e
	13'h0bd0: q2 = 16'h6f08; // 0x17a0
	13'h0bd1: q2 = 16'h3d7c; // 0x17a2
	13'h0bd2: q2 = 16'h0001; // 0x17a4
	13'h0bd3: q2 = 16'hffde; // 0x17a6
	13'h0bd4: q2 = 16'h6004; // 0x17a8
	13'h0bd5: q2 = 16'h426e; // 0x17aa
	13'h0bd6: q2 = 16'hffde; // 0x17ac
	13'h0bd7: q2 = 16'h4a6e; // 0x17ae
	13'h0bd8: q2 = 16'hffdc; // 0x17b0
	13'h0bd9: q2 = 16'h670a; // 0x17b2
	13'h0bda: q2 = 16'hbe7c; // 0x17b4
	13'h0bdb: q2 = 16'h0001; // 0x17b6
	13'h0bdc: q2 = 16'h6f04; // 0x17b8
	13'h0bdd: q2 = 16'h5347; // 0x17ba
	13'h0bde: q2 = 16'h6032; // 0x17bc
	13'h0bdf: q2 = 16'h4a6e; // 0x17be
	13'h0be0: q2 = 16'hffde; // 0x17c0
	13'h0be1: q2 = 16'h670a; // 0x17c2
	13'h0be2: q2 = 16'hbe6e; // 0x17c4
	13'h0be3: q2 = 16'hffe2; // 0x17c6
	13'h0be4: q2 = 16'h6c04; // 0x17c8
	13'h0be5: q2 = 16'h5247; // 0x17ca
	13'h0be6: q2 = 16'h6022; // 0x17cc
	13'h0be7: q2 = 16'h4a6e; // 0x17ce
	13'h0be8: q2 = 16'hffdc; // 0x17d0
	13'h0be9: q2 = 16'h670c; // 0x17d2
	13'h0bea: q2 = 16'hbc6e; // 0x17d4
	13'h0beb: q2 = 16'hfff8; // 0x17d6
	13'h0bec: q2 = 16'h6f06; // 0x17d8
	13'h0bed: q2 = 16'h536e; // 0x17da
	13'h0bee: q2 = 16'hfffe; // 0x17dc
	13'h0bef: q2 = 16'h6010; // 0x17de
	13'h0bf0: q2 = 16'h4a6e; // 0x17e0
	13'h0bf1: q2 = 16'hffde; // 0x17e2
	13'h0bf2: q2 = 16'h670a; // 0x17e4
	13'h0bf3: q2 = 16'hbc6e; // 0x17e6
	13'h0bf4: q2 = 16'hfff6; // 0x17e8
	13'h0bf5: q2 = 16'h6c04; // 0x17ea
	13'h0bf6: q2 = 16'h526e; // 0x17ec
	13'h0bf7: q2 = 16'hfffe; // 0x17ee
	13'h0bf8: q2 = 16'h4a79; // 0x17f0
	13'h0bf9: q2 = 16'h0001; // 0x17f2
	13'h0bfa: q2 = 16'h77e8; // 0x17f4
	13'h0bfb: q2 = 16'h6764; // 0x17f6
	13'h0bfc: q2 = 16'h2d79; // 0x17f8
	13'h0bfd: q2 = 16'h0000; // 0x17fa
	13'h0bfe: q2 = 16'hf96e; // 0x17fc
	13'h0bff: q2 = 16'hffd4; // 0x17fe
	13'h0c00: q2 = 16'h2039; // 0x1800
	13'h0c01: q2 = 16'h0000; // 0x1802
	13'h0c02: q2 = 16'hf972; // 0x1804
	13'h0c03: q2 = 16'he580; // 0x1806
	13'h0c04: q2 = 16'h91ae; // 0x1808
	13'h0c05: q2 = 16'hffd4; // 0x180a
	13'h0c06: q2 = 16'h206e; // 0x180c
	13'h0c07: q2 = 16'hffd4; // 0x180e
	13'h0c08: q2 = 16'h2010; // 0x1810
	13'h0c09: q2 = 16'h81fc; // 0x1812
	13'h0c0a: q2 = 16'h0e10; // 0x1814
	13'h0c0b: q2 = 16'h48c0; // 0x1816
	13'h0c0c: q2 = 16'hb0bc; // 0x1818
	13'h0c0d: q2 = 16'h0000; // 0x181a
	13'h0c0e: q2 = 16'h0014; // 0x181c
	13'h0c0f: q2 = 16'h663c; // 0x181e
	13'h0c10: q2 = 16'h206e; // 0x1820
	13'h0c11: q2 = 16'hffd4; // 0x1822
	13'h0c12: q2 = 16'h203c; // 0x1824
	13'h0c13: q2 = 16'h0000; // 0x1826
	13'h0c14: q2 = 16'h0e10; // 0x1828
	13'h0c15: q2 = 16'hd190; // 0x182a
	13'h0c16: q2 = 16'h2d7c; // 0x182c
	13'h0c17: q2 = 16'h0000; // 0x182e
	13'h0c18: q2 = 16'h7340; // 0x1830
	13'h0c19: q2 = 16'hffd8; // 0x1832
	13'h0c1a: q2 = 16'h2039; // 0x1834
	13'h0c1b: q2 = 16'h0000; // 0x1836
	13'h0c1c: q2 = 16'hf976; // 0x1838
	13'h0c1d: q2 = 16'he380; // 0x183a
	13'h0c1e: q2 = 16'hd1ae; // 0x183c
	13'h0c1f: q2 = 16'hffd8; // 0x183e
	13'h0c20: q2 = 16'h206e; // 0x1840
	13'h0c21: q2 = 16'hffd8; // 0x1842
	13'h0c22: q2 = 16'h30bc; // 0x1844
	13'h0c23: q2 = 16'h001b; // 0x1846
	13'h0c24: q2 = 16'h7017; // 0x1848
	13'h0c25: q2 = 16'h226e; // 0x184a
	13'h0c26: q2 = 16'hffd8; // 0x184c
	13'h0c27: q2 = 16'hd151; // 0x184e
	13'h0c28: q2 = 16'h206e; // 0x1850
	13'h0c29: q2 = 16'hffd8; // 0x1852
	13'h0c2a: q2 = 16'h226e; // 0x1854
	13'h0c2b: q2 = 16'hffd8; // 0x1856
	13'h0c2c: q2 = 16'h3151; // 0x1858
	13'h0c2d: q2 = 16'h0002; // 0x185a
	13'h0c2e: q2 = 16'h3c2e; // 0x185c
	13'h0c2f: q2 = 16'hfffe; // 0x185e
	13'h0c30: q2 = 16'hdc47; // 0x1860
	13'h0c31: q2 = 16'h5346; // 0x1862
	13'h0c32: q2 = 16'h302e; // 0x1864
	13'h0c33: q2 = 16'hfffe; // 0x1866
	13'h0c34: q2 = 16'hd07c; // 0x1868
	13'h0c35: q2 = 16'h000a; // 0x186a
	13'h0c36: q2 = 16'h5340; // 0x186c
	13'h0c37: q2 = 16'h3d40; // 0x186e
	13'h0c38: q2 = 16'hfffc; // 0x1870
	13'h0c39: q2 = 16'h4a6e; // 0x1872
	13'h0c3a: q2 = 16'hffdc; // 0x1874
	13'h0c3b: q2 = 16'h6712; // 0x1876
	13'h0c3c: q2 = 16'h4a44; // 0x1878
	13'h0c3d: q2 = 16'h6c04; // 0x187a
	13'h0c3e: q2 = 16'h5585; // 0x187c
	13'h0c3f: q2 = 16'h6006; // 0x187e
	13'h0c40: q2 = 16'h2a39; // 0x1880
	13'h0c41: q2 = 16'h0000; // 0x1882
	13'h0c42: q2 = 16'hf96a; // 0x1884
	13'h0c43: q2 = 16'h78ff; // 0x1886
	13'h0c44: q2 = 16'h6020; // 0x1888
	13'h0c45: q2 = 16'h4a6e; // 0x188a
	13'h0c46: q2 = 16'hffde; // 0x188c
	13'h0c47: q2 = 16'h6712; // 0x188e
	13'h0c48: q2 = 16'h4a44; // 0x1890
	13'h0c49: q2 = 16'h6f04; // 0x1892
	13'h0c4a: q2 = 16'h5585; // 0x1894
	13'h0c4b: q2 = 16'h6006; // 0x1896
	13'h0c4c: q2 = 16'h2a39; // 0x1898
	13'h0c4d: q2 = 16'h0000; // 0x189a
	13'h0c4e: q2 = 16'hf96a; // 0x189c
	13'h0c4f: q2 = 16'h7801; // 0x189e
	13'h0c50: q2 = 16'h6008; // 0x18a0
	13'h0c51: q2 = 16'h2a39; // 0x18a2
	13'h0c52: q2 = 16'h0000; // 0x18a4
	13'h0c53: q2 = 16'hf96a; // 0x18a6
	13'h0c54: q2 = 16'h4244; // 0x18a8
	13'h0c55: q2 = 16'h6000; // 0x18aa
	13'h0c56: q2 = 16'hfd9a; // 0x18ac
	13'h0c57: q2 = 16'h2079; // 0x18ae
	13'h0c58: q2 = 16'h0001; // 0x18b0
	13'h0c59: q2 = 16'h7fb8; // 0x18b2
	13'h0c5a: q2 = 16'h3086; // 0x18b4
	13'h0c5b: q2 = 16'h4a79; // 0x18b6
	13'h0c5c: q2 = 16'h0001; // 0x18b8
	13'h0c5d: q2 = 16'h7586; // 0x18ba
	13'h0c5e: q2 = 16'h673e; // 0x18bc
	13'h0c5f: q2 = 16'h2079; // 0x18be
	13'h0c60: q2 = 16'h0001; // 0x18c0
	13'h0c61: q2 = 16'h7fb8; // 0x18c2
	13'h0c62: q2 = 16'h3028; // 0x18c4
	13'h0c63: q2 = 16'h0002; // 0x18c6
	13'h0c64: q2 = 16'hb079; // 0x18c8
	13'h0c65: q2 = 16'h0001; // 0x18ca
	13'h0c66: q2 = 16'h7fce; // 0x18cc
	13'h0c67: q2 = 16'h6f2c; // 0x18ce
	13'h0c68: q2 = 16'h2079; // 0x18d0
	13'h0c69: q2 = 16'h0001; // 0x18d2
	13'h0c6a: q2 = 16'h7fb8; // 0x18d4
	13'h0c6b: q2 = 16'h3028; // 0x18d6
	13'h0c6c: q2 = 16'h0002; // 0x18d8
	13'h0c6d: q2 = 16'h9079; // 0x18da
	13'h0c6e: q2 = 16'h0001; // 0x18dc
	13'h0c6f: q2 = 16'h7fce; // 0x18de
	13'h0c70: q2 = 16'h48c0; // 0x18e0
	13'h0c71: q2 = 16'hd1b9; // 0x18e2
	13'h0c72: q2 = 16'h0001; // 0x18e4
	13'h0c73: q2 = 16'h75ba; // 0x18e6
	13'h0c74: q2 = 16'h3039; // 0x18e8
	13'h0c75: q2 = 16'h0001; // 0x18ea
	13'h0c76: q2 = 16'h8054; // 0x18ec
	13'h0c77: q2 = 16'he340; // 0x18ee
	13'h0c78: q2 = 16'h48c0; // 0x18f0
	13'h0c79: q2 = 16'hd0bc; // 0x18f2
	13'h0c7a: q2 = 16'h0001; // 0x18f4
	13'h0c7b: q2 = 16'h75da; // 0x18f6
	13'h0c7c: q2 = 16'h2040; // 0x18f8
	13'h0c7d: q2 = 16'h5250; // 0x18fa
	13'h0c7e: q2 = 16'h4eb9; // 0x18fc
	13'h0c7f: q2 = 16'h0000; // 0x18fe
	13'h0c80: q2 = 16'h0226; // 0x1900
	13'h0c81: q2 = 16'h4eb9; // 0x1902
	13'h0c82: q2 = 16'h0000; // 0x1904
	13'h0c83: q2 = 16'h8ea8; // 0x1906
	13'h0c84: q2 = 16'h4a9f; // 0x1908
	13'h0c85: q2 = 16'h4cdf; // 0x190a
	13'h0c86: q2 = 16'h00f8; // 0x190c
	13'h0c87: q2 = 16'h4e5e; // 0x190e
	13'h0c88: q2 = 16'h4e75; // 0x1910
	13'h0c89: q2 = 16'h4e56; // 0x1912
	13'h0c8a: q2 = 16'hfff2; // 0x1914
	13'h0c8b: q2 = 16'h48e7; // 0x1916
	13'h0c8c: q2 = 16'h0f04; // 0x1918
	13'h0c8d: q2 = 16'h4279; // 0x191a
	13'h0c8e: q2 = 16'h0001; // 0x191c
	13'h0c8f: q2 = 16'h7fc0; // 0x191e
	13'h0c90: q2 = 16'h2079; // 0x1920
	13'h0c91: q2 = 16'h0001; // 0x1922
	13'h0c92: q2 = 16'h7fb8; // 0x1924
	13'h0c93: q2 = 16'h33e8; // 0x1926
	13'h0c94: q2 = 16'h0002; // 0x1928
	13'h0c95: q2 = 16'h0001; // 0x192a
	13'h0c96: q2 = 16'h7fce; // 0x192c
	13'h0c97: q2 = 16'h7e01; // 0x192e
	13'h0c98: q2 = 16'h3d7c; // 0x1930
	13'h0c99: q2 = 16'h0034; // 0x1932
	13'h0c9a: q2 = 16'hfffc; // 0x1934
	13'h0c9b: q2 = 16'hbe7c; // 0x1936
	13'h0c9c: q2 = 16'h000a; // 0x1938
	13'h0c9d: q2 = 16'h6e2c; // 0x193a
	13'h0c9e: q2 = 16'h3eae; // 0x193c
	13'h0c9f: q2 = 16'hfffc; // 0x193e
	13'h0ca0: q2 = 16'h200e; // 0x1940
	13'h0ca1: q2 = 16'hd0bc; // 0x1942
	13'h0ca2: q2 = 16'hffff; // 0x1944
	13'h0ca3: q2 = 16'hfff2; // 0x1946
	13'h0ca4: q2 = 16'h2f00; // 0x1948
	13'h0ca5: q2 = 16'h200e; // 0x194a
	13'h0ca6: q2 = 16'hd0bc; // 0x194c
	13'h0ca7: q2 = 16'hffff; // 0x194e
	13'h0ca8: q2 = 16'hfff8; // 0x1950
	13'h0ca9: q2 = 16'h2f00; // 0x1952
	13'h0caa: q2 = 16'h3f07; // 0x1954
	13'h0cab: q2 = 16'h4eb9; // 0x1956
	13'h0cac: q2 = 16'h0000; // 0x1958
	13'h0cad: q2 = 16'h1402; // 0x195a
	13'h0cae: q2 = 16'hdefc; // 0x195c
	13'h0caf: q2 = 16'h000a; // 0x195e
	13'h0cb0: q2 = 16'h5247; // 0x1960
	13'h0cb1: q2 = 16'h526e; // 0x1962
	13'h0cb2: q2 = 16'hfffc; // 0x1964
	13'h0cb3: q2 = 16'h60ce; // 0x1966
	13'h0cb4: q2 = 16'h2a7c; // 0x1968
	13'h0cb5: q2 = 16'h0000; // 0x196a
	13'h0cb6: q2 = 16'hf97c; // 0x196c
	13'h0cb7: q2 = 16'h7c12; // 0x196e
	13'h0cb8: q2 = 16'hbc7c; // 0x1970
	13'h0cb9: q2 = 16'h000c; // 0x1972
	13'h0cba: q2 = 16'h6d3c; // 0x1974
	13'h0cbb: q2 = 16'h7e04; // 0x1976
	13'h0cbc: q2 = 16'hbe7c; // 0x1978
	13'h0cbd: q2 = 16'h000a; // 0x197a
	13'h0cbe: q2 = 16'h6e30; // 0x197c
	13'h0cbf: q2 = 16'h1015; // 0x197e
	13'h0cc0: q2 = 16'h4880; // 0x1980
	13'h0cc1: q2 = 16'h3d40; // 0x1982
	13'h0cc2: q2 = 16'hfffe; // 0x1984
	13'h0cc3: q2 = 16'h0c6e; // 0x1986
	13'h0cc4: q2 = 16'h0020; // 0x1988
	13'h0cc5: q2 = 16'hfffe; // 0x198a
	13'h0cc6: q2 = 16'h6c06; // 0x198c
	13'h0cc7: q2 = 16'h066e; // 0x198e
	13'h0cc8: q2 = 16'h0100; // 0x1990
	13'h0cc9: q2 = 16'hfffe; // 0x1992
	13'h0cca: q2 = 16'h3ebc; // 0x1994
	13'h0ccb: q2 = 16'h0021; // 0x1996
	13'h0ccc: q2 = 16'h3f2e; // 0x1998
	13'h0ccd: q2 = 16'hfffe; // 0x199a
	13'h0cce: q2 = 16'h3f06; // 0x199c
	13'h0ccf: q2 = 16'h3f07; // 0x199e
	13'h0cd0: q2 = 16'h4eb9; // 0x19a0
	13'h0cd1: q2 = 16'h0000; // 0x19a2
	13'h0cd2: q2 = 16'h3d18; // 0x19a4
	13'h0cd3: q2 = 16'h5c4f; // 0x19a6
	13'h0cd4: q2 = 16'h5247; // 0x19a8
	13'h0cd5: q2 = 16'h528d; // 0x19aa
	13'h0cd6: q2 = 16'h60ca; // 0x19ac
	13'h0cd7: q2 = 16'h5346; // 0x19ae
	13'h0cd8: q2 = 16'h60be; // 0x19b0
	13'h0cd9: q2 = 16'h3d7c; // 0x19b2
	13'h0cda: q2 = 16'h0002; // 0x19b4
	13'h0cdb: q2 = 16'hfffa; // 0x19b6
	13'h0cdc: q2 = 16'h3a2e; // 0x19b8
	13'h0cdd: q2 = 16'hfffa; // 0x19ba
	13'h0cde: q2 = 16'h4247; // 0x19bc
	13'h0cdf: q2 = 16'hbe7c; // 0x19be
	13'h0ce0: q2 = 16'h000a; // 0x19c0
	13'h0ce1: q2 = 16'h6c1c; // 0x19c2
	13'h0ce2: q2 = 16'h3ebc; // 0x19c4
	13'h0ce3: q2 = 16'h0021; // 0x19c6
	13'h0ce4: q2 = 16'h3f3c; // 0x19c8
	13'h0ce5: q2 = 16'h00d8; // 0x19ca
	13'h0ce6: q2 = 16'h3f3c; // 0x19cc
	13'h0ce7: q2 = 16'h0009; // 0x19ce
	13'h0ce8: q2 = 16'h3f05; // 0x19d0
	13'h0ce9: q2 = 16'h4eb9; // 0x19d2
	13'h0cea: q2 = 16'h0000; // 0x19d4
	13'h0ceb: q2 = 16'h3d18; // 0x19d6
	13'h0cec: q2 = 16'h5c4f; // 0x19d8
	13'h0ced: q2 = 16'h5645; // 0x19da
	13'h0cee: q2 = 16'h5247; // 0x19dc
	13'h0cef: q2 = 16'h60de; // 0x19de
	13'h0cf0: q2 = 16'h7e01; // 0x19e0
	13'h0cf1: q2 = 16'hbe7c; // 0x19e2
	13'h0cf2: q2 = 16'h0003; // 0x19e4
	13'h0cf3: q2 = 16'h6e0c; // 0x19e6
	13'h0cf4: q2 = 16'h3e87; // 0x19e8
	13'h0cf5: q2 = 16'h4eb9; // 0x19ea
	13'h0cf6: q2 = 16'h0000; // 0x19ec
	13'h0cf7: q2 = 16'h8a22; // 0x19ee
	13'h0cf8: q2 = 16'h5247; // 0x19f0
	13'h0cf9: q2 = 16'h60ee; // 0x19f2
	13'h0cfa: q2 = 16'h4a9f; // 0x19f4
	13'h0cfb: q2 = 16'h4cdf; // 0x19f6
	13'h0cfc: q2 = 16'h20e0; // 0x19f8
	13'h0cfd: q2 = 16'h4e5e; // 0x19fa
	13'h0cfe: q2 = 16'h4e75; // 0x19fc
	13'h0cff: q2 = 16'h4e56; // 0x19fe
	13'h0d00: q2 = 16'h0000; // 0x1a00
	13'h0d01: q2 = 16'h48e7; // 0x1a02
	13'h0d02: q2 = 16'h1f00; // 0x1a04
	13'h0d03: q2 = 16'h4279; // 0x1a06
	13'h0d04: q2 = 16'h0001; // 0x1a08
	13'h0d05: q2 = 16'h76d6; // 0x1a0a
	13'h0d06: q2 = 16'h7c04; // 0x1a0c
	13'h0d07: q2 = 16'hbc7c; // 0x1a0e
	13'h0d08: q2 = 16'h001f; // 0x1a10
	13'h0d09: q2 = 16'h6e24; // 0x1a12
	13'h0d0a: q2 = 16'h4247; // 0x1a14
	13'h0d0b: q2 = 16'hbe7c; // 0x1a16
	13'h0d0c: q2 = 16'h001f; // 0x1a18
	13'h0d0d: q2 = 16'h6e18; // 0x1a1a
	13'h0d0e: q2 = 16'h3ebc; // 0x1a1c
	13'h0d0f: q2 = 16'h001d; // 0x1a1e
	13'h0d10: q2 = 16'h3f3c; // 0x1a20
	13'h0d11: q2 = 16'h0003; // 0x1a22
	13'h0d12: q2 = 16'h3f06; // 0x1a24
	13'h0d13: q2 = 16'h3f07; // 0x1a26
	13'h0d14: q2 = 16'h4eb9; // 0x1a28
	13'h0d15: q2 = 16'h0000; // 0x1a2a
	13'h0d16: q2 = 16'h3d18; // 0x1a2c
	13'h0d17: q2 = 16'h5c4f; // 0x1a2e
	13'h0d18: q2 = 16'h5247; // 0x1a30
	13'h0d19: q2 = 16'h60e2; // 0x1a32
	13'h0d1a: q2 = 16'h5246; // 0x1a34
	13'h0d1b: q2 = 16'h60d6; // 0x1a36
	13'h0d1c: q2 = 16'h4244; // 0x1a38
	13'h0d1d: q2 = 16'h7c08; // 0x1a3a
	13'h0d1e: q2 = 16'hbc7c; // 0x1a3c
	13'h0d1f: q2 = 16'h0018; // 0x1a3e
	13'h0d20: q2 = 16'h6c00; // 0x1a40
	13'h0d21: q2 = 16'h007e; // 0x1a42
	13'h0d22: q2 = 16'h7e08; // 0x1a44
	13'h0d23: q2 = 16'hbe7c; // 0x1a46
	13'h0d24: q2 = 16'h0018; // 0x1a48
	13'h0d25: q2 = 16'h6c6e; // 0x1a4a
	13'h0d26: q2 = 16'h3007; // 0x1a4c
	13'h0d27: q2 = 16'hc07c; // 0x1a4e
	13'h0d28: q2 = 16'h0010; // 0x1a50
	13'h0d29: q2 = 16'he540; // 0x1a52
	13'h0d2a: q2 = 16'h3206; // 0x1a54
	13'h0d2b: q2 = 16'hc27c; // 0x1a56
	13'h0d2c: q2 = 16'h0010; // 0x1a58
	13'h0d2d: q2 = 16'he741; // 0x1a5a
	13'h0d2e: q2 = 16'h8041; // 0x1a5c
	13'h0d2f: q2 = 16'h3a00; // 0x1a5e
	13'h0d30: q2 = 16'hbc7c; // 0x1a60
	13'h0d31: q2 = 16'h0010; // 0x1a62
	13'h0d32: q2 = 16'h6c06; // 0x1a64
	13'h0d33: q2 = 16'h700f; // 0x1a66
	13'h0d34: q2 = 16'h9046; // 0x1a68
	13'h0d35: q2 = 16'h6006; // 0x1a6a
	13'h0d36: q2 = 16'h3006; // 0x1a6c
	13'h0d37: q2 = 16'hd07c; // 0x1a6e
	13'h0d38: q2 = 16'hfff0; // 0x1a70
	13'h0d39: q2 = 16'he740; // 0x1a72
	13'h0d3a: q2 = 16'h8a40; // 0x1a74
	13'h0d3b: q2 = 16'hbe7c; // 0x1a76
	13'h0d3c: q2 = 16'h0010; // 0x1a78
	13'h0d3d: q2 = 16'h6c06; // 0x1a7a
	13'h0d3e: q2 = 16'h700f; // 0x1a7c
	13'h0d3f: q2 = 16'h9047; // 0x1a7e
	13'h0d40: q2 = 16'h6006; // 0x1a80
	13'h0d41: q2 = 16'h3007; // 0x1a82
	13'h0d42: q2 = 16'hd07c; // 0x1a84
	13'h0d43: q2 = 16'hfff0; // 0x1a86
	13'h0d44: q2 = 16'h8a40; // 0x1a88
	13'h0d45: q2 = 16'h3004; // 0x1a8a
	13'h0d46: q2 = 16'he340; // 0x1a8c
	13'h0d47: q2 = 16'h48c0; // 0x1a8e
	13'h0d48: q2 = 16'hd0bc; // 0x1a90
	13'h0d49: q2 = 16'h0001; // 0x1a92
	13'h0d4a: q2 = 16'h75e8; // 0x1a94
	13'h0d4b: q2 = 16'h2040; // 0x1a96
	13'h0d4c: q2 = 16'h3085; // 0x1a98
	13'h0d4d: q2 = 16'h3004; // 0x1a9a
	13'h0d4e: q2 = 16'he440; // 0x1a9c
	13'h0d4f: q2 = 16'h3e80; // 0x1a9e
	13'h0d50: q2 = 16'h3f07; // 0x1aa0
	13'h0d51: q2 = 16'h0257; // 0x1aa2
	13'h0d52: q2 = 16'h0003; // 0x1aa4
	13'h0d53: q2 = 16'h3f06; // 0x1aa6
	13'h0d54: q2 = 16'h5457; // 0x1aa8
	13'h0d55: q2 = 16'h3f07; // 0x1aaa
	13'h0d56: q2 = 16'h4eb9; // 0x1aac
	13'h0d57: q2 = 16'h0000; // 0x1aae
	13'h0d58: q2 = 16'h3d18; // 0x1ab0
	13'h0d59: q2 = 16'h5c4f; // 0x1ab2
	13'h0d5a: q2 = 16'h5244; // 0x1ab4
	13'h0d5b: q2 = 16'h5247; // 0x1ab6
	13'h0d5c: q2 = 16'h608c; // 0x1ab8
	13'h0d5d: q2 = 16'h5246; // 0x1aba
	13'h0d5e: q2 = 16'h6000; // 0x1abc
	13'h0d5f: q2 = 16'hff7e; // 0x1abe
	13'h0d60: q2 = 16'h4a79; // 0x1ac0
	13'h0d61: q2 = 16'h0001; // 0x1ac2
	13'h0d62: q2 = 16'h8a7e; // 0x1ac4
	13'h0d63: q2 = 16'h6702; // 0x1ac6
	13'h0d64: q2 = 16'h60f6; // 0x1ac8
	13'h0d65: q2 = 16'h4a79; // 0x1aca
	13'h0d66: q2 = 16'h0001; // 0x1acc
	13'h0d67: q2 = 16'h8a7e; // 0x1ace
	13'h0d68: q2 = 16'h6602; // 0x1ad0
	13'h0d69: q2 = 16'h60f6; // 0x1ad2
	13'h0d6a: q2 = 16'h4eb9; // 0x1ad4
	13'h0d6b: q2 = 16'h0000; // 0x1ad6
	13'h0d6c: q2 = 16'h8ea8; // 0x1ad8
	13'h0d6d: q2 = 16'h4a9f; // 0x1ada
	13'h0d6e: q2 = 16'h4cdf; // 0x1adc
	13'h0d6f: q2 = 16'h00f0; // 0x1ade
	13'h0d70: q2 = 16'h4e5e; // 0x1ae0
	13'h0d71: q2 = 16'h4e75; // 0x1ae2
	13'h0d72: q2 = 16'h4e56; // 0x1ae4
	13'h0d73: q2 = 16'h0000; // 0x1ae6
	13'h0d74: q2 = 16'h48e7; // 0x1ae8
	13'h0d75: q2 = 16'h0f00; // 0x1aea
	13'h0d76: q2 = 16'h7c04; // 0x1aec
	13'h0d77: q2 = 16'hbc7c; // 0x1aee
	13'h0d78: q2 = 16'h001f; // 0x1af0
	13'h0d79: q2 = 16'h6e3e; // 0x1af2
	13'h0d7a: q2 = 16'h4247; // 0x1af4
	13'h0d7b: q2 = 16'hbe7c; // 0x1af6
	13'h0d7c: q2 = 16'h001f; // 0x1af8
	13'h0d7d: q2 = 16'h6e32; // 0x1afa
	13'h0d7e: q2 = 16'h7a0c; // 0x1afc
	13'h0d7f: q2 = 16'h3006; // 0x1afe
	13'h0d80: q2 = 16'hc07c; // 0x1b00
	13'h0d81: q2 = 16'h0001; // 0x1b02
	13'h0d82: q2 = 16'h7201; // 0x1b04
	13'h0d83: q2 = 16'hb340; // 0x1b06
	13'h0d84: q2 = 16'h8a40; // 0x1b08
	13'h0d85: q2 = 16'h3007; // 0x1b0a
	13'h0d86: q2 = 16'hc07c; // 0x1b0c
	13'h0d87: q2 = 16'h0001; // 0x1b0e
	13'h0d88: q2 = 16'h7201; // 0x1b10
	13'h0d89: q2 = 16'hb340; // 0x1b12
	13'h0d8a: q2 = 16'he340; // 0x1b14
	13'h0d8b: q2 = 16'h8a40; // 0x1b16
	13'h0d8c: q2 = 16'h3ebc; // 0x1b18
	13'h0d8d: q2 = 16'h003e; // 0x1b1a
	13'h0d8e: q2 = 16'h3f05; // 0x1b1c
	13'h0d8f: q2 = 16'h3f06; // 0x1b1e
	13'h0d90: q2 = 16'h3f07; // 0x1b20
	13'h0d91: q2 = 16'h4eb9; // 0x1b22
	13'h0d92: q2 = 16'h0000; // 0x1b24
	13'h0d93: q2 = 16'h3d18; // 0x1b26
	13'h0d94: q2 = 16'h5c4f; // 0x1b28
	13'h0d95: q2 = 16'h5247; // 0x1b2a
	13'h0d96: q2 = 16'h60c8; // 0x1b2c
	13'h0d97: q2 = 16'h5246; // 0x1b2e
	13'h0d98: q2 = 16'h60bc; // 0x1b30
	13'h0d99: q2 = 16'h4a79; // 0x1b32
	13'h0d9a: q2 = 16'h0001; // 0x1b34
	13'h0d9b: q2 = 16'h8a7e; // 0x1b36
	13'h0d9c: q2 = 16'h6702; // 0x1b38
	13'h0d9d: q2 = 16'h60f6; // 0x1b3a
	13'h0d9e: q2 = 16'h4a79; // 0x1b3c
	13'h0d9f: q2 = 16'h0001; // 0x1b3e
	13'h0da0: q2 = 16'h8a7e; // 0x1b40
	13'h0da1: q2 = 16'h6602; // 0x1b42
	13'h0da2: q2 = 16'h60f6; // 0x1b44
	13'h0da3: q2 = 16'h4a9f; // 0x1b46
	13'h0da4: q2 = 16'h4cdf; // 0x1b48
	13'h0da5: q2 = 16'h00e0; // 0x1b4a
	13'h0da6: q2 = 16'h4e5e; // 0x1b4c
	13'h0da7: q2 = 16'h4e75; // 0x1b4e
	13'h0da8: q2 = 16'h4e56; // 0x1b50
	13'h0da9: q2 = 16'hffde; // 0x1b52
	13'h0daa: q2 = 16'h48e7; // 0x1b54
	13'h0dab: q2 = 16'h1f04; // 0x1b56
	13'h0dac: q2 = 16'h4eb9; // 0x1b58
	13'h0dad: q2 = 16'h0000; // 0x1b5a
	13'h0dae: q2 = 16'h0226; // 0x1b5c
	13'h0daf: q2 = 16'h7801; // 0x1b5e
	13'h0db0: q2 = 16'h4247; // 0x1b60
	13'h0db1: q2 = 16'hbe7c; // 0x1b62
	13'h0db2: q2 = 16'h0005; // 0x1b64
	13'h0db3: q2 = 16'h6e62; // 0x1b66
	13'h0db4: q2 = 16'h4a79; // 0x1b68
	13'h0db5: q2 = 16'h0001; // 0x1b6a
	13'h0db6: q2 = 16'h758e; // 0x1b6c
	13'h0db7: q2 = 16'h660c; // 0x1b6e
	13'h0db8: q2 = 16'hbe7c; // 0x1b70
	13'h0db9: q2 = 16'h0003; // 0x1b72
	13'h0dba: q2 = 16'h6750; // 0x1b74
	13'h0dbb: q2 = 16'hbe7c; // 0x1b76
	13'h0dbc: q2 = 16'h0004; // 0x1b78
	13'h0dbd: q2 = 16'h674a; // 0x1b7a
	13'h0dbe: q2 = 16'h3eb9; // 0x1b7c
	13'h0dbf: q2 = 16'h0000; // 0x1b7e
	13'h0dc0: q2 = 16'hf9ce; // 0x1b80
	13'h0dc1: q2 = 16'h3007; // 0x1b82
	13'h0dc2: q2 = 16'hd157; // 0x1b84
	13'h0dc3: q2 = 16'h200e; // 0x1b86
	13'h0dc4: q2 = 16'hd0bc; // 0x1b88
	13'h0dc5: q2 = 16'hffff; // 0x1b8a
	13'h0dc6: q2 = 16'hffde; // 0x1b8c
	13'h0dc7: q2 = 16'h2f00; // 0x1b8e
	13'h0dc8: q2 = 16'h4eb9; // 0x1b90
	13'h0dc9: q2 = 16'h0000; // 0x1b92
	13'h0dca: q2 = 16'h78f6; // 0x1b94
	13'h0dcb: q2 = 16'h4a9f; // 0x1b96
	13'h0dcc: q2 = 16'h3ebc; // 0x1b98
	13'h0dcd: q2 = 16'h0036; // 0x1b9a
	13'h0dce: q2 = 16'h4267; // 0x1b9c
	13'h0dcf: q2 = 16'h3f3c; // 0x1b9e
	13'h0dd0: q2 = 16'h0064; // 0x1ba0
	13'h0dd1: q2 = 16'h3007; // 0x1ba2
	13'h0dd2: q2 = 16'he340; // 0x1ba4
	13'h0dd3: q2 = 16'h48c0; // 0x1ba6
	13'h0dd4: q2 = 16'hd0bc; // 0x1ba8
	13'h0dd5: q2 = 16'h0000; // 0x1baa
	13'h0dd6: q2 = 16'hf9d0; // 0x1bac
	13'h0dd7: q2 = 16'h2040; // 0x1bae
	13'h0dd8: q2 = 16'h3f10; // 0x1bb0
	13'h0dd9: q2 = 16'h200e; // 0x1bb2
	13'h0dda: q2 = 16'hd0bc; // 0x1bb4
	13'h0ddb: q2 = 16'hffff; // 0x1bb6
	13'h0ddc: q2 = 16'hffde; // 0x1bb8
	13'h0ddd: q2 = 16'h2f00; // 0x1bba
	13'h0dde: q2 = 16'h4eb9; // 0x1bbc
	13'h0ddf: q2 = 16'h0000; // 0x1bbe
	13'h0de0: q2 = 16'h026c; // 0x1bc0
	13'h0de1: q2 = 16'hdefc; // 0x1bc2
	13'h0de2: q2 = 16'h000a; // 0x1bc4
	13'h0de3: q2 = 16'h5247; // 0x1bc6
	13'h0de4: q2 = 16'h6098; // 0x1bc8
	13'h0de5: q2 = 16'h4a79; // 0x1bca
	13'h0de6: q2 = 16'h0001; // 0x1bcc
	13'h0de7: q2 = 16'h758e; // 0x1bce
	13'h0de8: q2 = 16'h6718; // 0x1bd0
	13'h0de9: q2 = 16'h3ebc; // 0x1bd2
	13'h0dea: q2 = 16'h0036; // 0x1bd4
	13'h0deb: q2 = 16'h3f3c; // 0x1bd6
	13'h0dec: q2 = 16'h0032; // 0x1bd8
	13'h0ded: q2 = 16'h3f3c; // 0x1bda
	13'h0dee: q2 = 16'h0010; // 0x1bdc
	13'h0def: q2 = 16'h3f3c; // 0x1bde
	13'h0df0: q2 = 16'h000f; // 0x1be0
	13'h0df1: q2 = 16'h4eb9; // 0x1be2
	13'h0df2: q2 = 16'h0000; // 0x1be4
	13'h0df3: q2 = 16'h3d18; // 0x1be6
	13'h0df4: q2 = 16'h5c4f; // 0x1be8
	13'h0df5: q2 = 16'h7c01; // 0x1bea
	13'h0df6: q2 = 16'h7a01; // 0x1bec
	13'h0df7: q2 = 16'h2a7c; // 0x1bee
	13'h0df8: q2 = 16'h0001; // 0x1bf0
	13'h0df9: q2 = 16'h8684; // 0x1bf2
	13'h0dfa: q2 = 16'h4247; // 0x1bf4
	13'h0dfb: q2 = 16'hbe7c; // 0x1bf6
	13'h0dfc: q2 = 16'h0008; // 0x1bf8
	13'h0dfd: q2 = 16'h6c0a; // 0x1bfa
	13'h0dfe: q2 = 16'h3abc; // 0x1bfc
	13'h0dff: q2 = 16'h0080; // 0x1bfe
	13'h0e00: q2 = 16'h5247; // 0x1c00
	13'h0e01: q2 = 16'h548d; // 0x1c02
	13'h0e02: q2 = 16'h60f0; // 0x1c04
	13'h0e03: q2 = 16'h4240; // 0x1c06
	13'h0e04: q2 = 16'h33c0; // 0x1c08
	13'h0e05: q2 = 16'h0001; // 0x1c0a
	13'h0e06: q2 = 16'h86aa; // 0x1c0c
	13'h0e07: q2 = 16'h33c0; // 0x1c0e
	13'h0e08: q2 = 16'h0001; // 0x1c10
	13'h0e09: q2 = 16'h8680; // 0x1c12
	13'h0e0a: q2 = 16'h4a46; // 0x1c14
	13'h0e0b: q2 = 16'h6608; // 0x1c16
	13'h0e0c: q2 = 16'h4a79; // 0x1c18
	13'h0e0d: q2 = 16'h0001; // 0x1c1a
	13'h0e0e: q2 = 16'h8a7e; // 0x1c1c
	13'h0e0f: q2 = 16'h665a; // 0x1c1e
	13'h0e10: q2 = 16'h4a45; // 0x1c20
	13'h0e11: q2 = 16'h6640; // 0x1c22
	13'h0e12: q2 = 16'h4a79; // 0x1c24
	13'h0e13: q2 = 16'h0001; // 0x1c26
	13'h0e14: q2 = 16'h8a80; // 0x1c28
	13'h0e15: q2 = 16'h6738; // 0x1c2a
	13'h0e16: q2 = 16'h4a79; // 0x1c2c
	13'h0e17: q2 = 16'h0001; // 0x1c2e
	13'h0e18: q2 = 16'h758e; // 0x1c30
	13'h0e19: q2 = 16'h6730; // 0x1c32
	13'h0e1a: q2 = 16'h7001; // 0x1c34
	13'h0e1b: q2 = 16'h9079; // 0x1c36
	13'h0e1c: q2 = 16'h0001; // 0x1c38
	13'h0e1d: q2 = 16'h8052; // 0x1c3a
	13'h0e1e: q2 = 16'h33c0; // 0x1c3c
	13'h0e1f: q2 = 16'h0001; // 0x1c3e
	13'h0e20: q2 = 16'h8052; // 0x1c40
	13'h0e21: q2 = 16'h7001; // 0x1c42
	13'h0e22: q2 = 16'h9044; // 0x1c44
	13'h0e23: q2 = 16'h3800; // 0x1c46
	13'h0e24: q2 = 16'h7a01; // 0x1c48
	13'h0e25: q2 = 16'h3ebc; // 0x1c4a
	13'h0e26: q2 = 16'h0036; // 0x1c4c
	13'h0e27: q2 = 16'h3f04; // 0x1c4e
	13'h0e28: q2 = 16'h0657; // 0x1c50
	13'h0e29: q2 = 16'h0031; // 0x1c52
	13'h0e2a: q2 = 16'h3f3c; // 0x1c54
	13'h0e2b: q2 = 16'h0010; // 0x1c56
	13'h0e2c: q2 = 16'h3f3c; // 0x1c58
	13'h0e2d: q2 = 16'h000f; // 0x1c5a
	13'h0e2e: q2 = 16'h4eb9; // 0x1c5c
	13'h0e2f: q2 = 16'h0000; // 0x1c5e
	13'h0e30: q2 = 16'h3d18; // 0x1c60
	13'h0e31: q2 = 16'h5c4f; // 0x1c62
	13'h0e32: q2 = 16'h4a79; // 0x1c64
	13'h0e33: q2 = 16'h0001; // 0x1c66
	13'h0e34: q2 = 16'h8a7e; // 0x1c68
	13'h0e35: q2 = 16'h6602; // 0x1c6a
	13'h0e36: q2 = 16'h4246; // 0x1c6c
	13'h0e37: q2 = 16'h4a79; // 0x1c6e
	13'h0e38: q2 = 16'h0001; // 0x1c70
	13'h0e39: q2 = 16'h8a80; // 0x1c72
	13'h0e3a: q2 = 16'h6602; // 0x1c74
	13'h0e3b: q2 = 16'h4245; // 0x1c76
	13'h0e3c: q2 = 16'h609a; // 0x1c78
	13'h0e3d: q2 = 16'h4279; // 0x1c7a
	13'h0e3e: q2 = 16'h0001; // 0x1c7c
	13'h0e3f: q2 = 16'h8052; // 0x1c7e
	13'h0e40: q2 = 16'h4a9f; // 0x1c80
	13'h0e41: q2 = 16'h4cdf; // 0x1c82
	13'h0e42: q2 = 16'h20f0; // 0x1c84
	13'h0e43: q2 = 16'h4e5e; // 0x1c86
	13'h0e44: q2 = 16'h4e75; // 0x1c88
	13'h0e45: q2 = 16'h4e56; // 0x1c8a
	13'h0e46: q2 = 16'hffde; // 0x1c8c
	13'h0e47: q2 = 16'h48e7; // 0x1c8e
	13'h0e48: q2 = 16'h3f00; // 0x1c90
	13'h0e49: q2 = 16'h4eb9; // 0x1c92
	13'h0e4a: q2 = 16'h0000; // 0x1c94
	13'h0e4b: q2 = 16'h0226; // 0x1c96
	13'h0e4c: q2 = 16'h4eb9; // 0x1c98
	13'h0e4d: q2 = 16'h0000; // 0x1c9a
	13'h0e4e: q2 = 16'h8ea8; // 0x1c9c
	13'h0e4f: q2 = 16'h4eb9; // 0x1c9e
	13'h0e50: q2 = 16'h0000; // 0x1ca0
	13'h0e51: q2 = 16'had94; // 0x1ca2
	13'h0e52: q2 = 16'h4eb9; // 0x1ca4
	13'h0e53: q2 = 16'h0000; // 0x1ca6
	13'h0e54: q2 = 16'had94; // 0x1ca8
	13'h0e55: q2 = 16'h4eb9; // 0x1caa
	13'h0e56: q2 = 16'h0000; // 0x1cac
	13'h0e57: q2 = 16'h8902; // 0x1cae
	13'h0e58: q2 = 16'h33fc; // 0x1cb0
	13'h0e59: q2 = 16'h0001; // 0x1cb2
	13'h0e5a: q2 = 16'h0001; // 0x1cb4
	13'h0e5b: q2 = 16'h8a7a; // 0x1cb6
	13'h0e5c: q2 = 16'h4279; // 0x1cb8
	13'h0e5d: q2 = 16'h0001; // 0x1cba
	13'h0e5e: q2 = 16'h7fa6; // 0x1cbc
	13'h0e5f: q2 = 16'h4279; // 0x1cbe
	13'h0e60: q2 = 16'h0001; // 0x1cc0
	13'h0e61: q2 = 16'h8052; // 0x1cc2
	13'h0e62: q2 = 16'h33fc; // 0x1cc4
	13'h0e63: q2 = 16'h0001; // 0x1cc6
	13'h0e64: q2 = 16'h0001; // 0x1cc8
	13'h0e65: q2 = 16'h85fc; // 0x1cca
	13'h0e66: q2 = 16'h4246; // 0x1ccc
	13'h0e67: q2 = 16'h7a01; // 0x1cce
	13'h0e68: q2 = 16'h4247; // 0x1cd0
	13'h0e69: q2 = 16'hbe7c; // 0x1cd2
	13'h0e6a: q2 = 16'h0006; // 0x1cd4
	13'h0e6b: q2 = 16'h6e60; // 0x1cd6
	13'h0e6c: q2 = 16'hbe46; // 0x1cd8
	13'h0e6d: q2 = 16'h6604; // 0x1cda
	13'h0e6e: q2 = 16'h782d; // 0x1cdc
	13'h0e6f: q2 = 16'h6002; // 0x1cde
	13'h0e70: q2 = 16'h7836; // 0x1ce0
	13'h0e71: q2 = 16'hbe7c; // 0x1ce2
	13'h0e72: q2 = 16'h0002; // 0x1ce4
	13'h0e73: q2 = 16'h6e04; // 0x1ce6
	13'h0e74: q2 = 16'h760c; // 0x1ce8
	13'h0e75: q2 = 16'h6002; // 0x1cea
	13'h0e76: q2 = 16'h7664; // 0x1cec
	13'h0e77: q2 = 16'h3eb9; // 0x1cee
	13'h0e78: q2 = 16'h0000; // 0x1cf0
	13'h0e79: q2 = 16'hf9ae; // 0x1cf2
	13'h0e7a: q2 = 16'h3007; // 0x1cf4
	13'h0e7b: q2 = 16'hd157; // 0x1cf6
	13'h0e7c: q2 = 16'h200e; // 0x1cf8
	13'h0e7d: q2 = 16'hd0bc; // 0x1cfa
	13'h0e7e: q2 = 16'hffff; // 0x1cfc
	13'h0e7f: q2 = 16'hffde; // 0x1cfe
	13'h0e80: q2 = 16'h2f00; // 0x1d00
	13'h0e81: q2 = 16'h4eb9; // 0x1d02
	13'h0e82: q2 = 16'h0000; // 0x1d04
	13'h0e83: q2 = 16'h78f6; // 0x1d06
	13'h0e84: q2 = 16'h4a9f; // 0x1d08
	13'h0e85: q2 = 16'h3e84; // 0x1d0a
	13'h0e86: q2 = 16'h4267; // 0x1d0c
	13'h0e87: q2 = 16'h3f03; // 0x1d0e
	13'h0e88: q2 = 16'h3007; // 0x1d10
	13'h0e89: q2 = 16'he340; // 0x1d12
	13'h0e8a: q2 = 16'h48c0; // 0x1d14
	13'h0e8b: q2 = 16'hd0bc; // 0x1d16
	13'h0e8c: q2 = 16'h0000; // 0x1d18
	13'h0e8d: q2 = 16'hf9b0; // 0x1d1a
	13'h0e8e: q2 = 16'h2040; // 0x1d1c
	13'h0e8f: q2 = 16'h3f10; // 0x1d1e
	13'h0e90: q2 = 16'h200e; // 0x1d20
	13'h0e91: q2 = 16'hd0bc; // 0x1d22
	13'h0e92: q2 = 16'hffff; // 0x1d24
	13'h0e93: q2 = 16'hffde; // 0x1d26
	13'h0e94: q2 = 16'h2f00; // 0x1d28
	13'h0e95: q2 = 16'h4eb9; // 0x1d2a
	13'h0e96: q2 = 16'h0000; // 0x1d2c
	13'h0e97: q2 = 16'h026c; // 0x1d2e
	13'h0e98: q2 = 16'hdefc; // 0x1d30
	13'h0e99: q2 = 16'h000a; // 0x1d32
	13'h0e9a: q2 = 16'h5247; // 0x1d34
	13'h0e9b: q2 = 16'h609a; // 0x1d36
	13'h0e9c: q2 = 16'h3ebc; // 0x1d38
	13'h0e9d: q2 = 16'h0002; // 0x1d3a
	13'h0e9e: q2 = 16'h3f06; // 0x1d3c
	13'h0e9f: q2 = 16'h4eb9; // 0x1d3e
	13'h0ea0: q2 = 16'h0000; // 0x1d40
	13'h0ea1: q2 = 16'ha602; // 0x1d42
	13'h0ea2: q2 = 16'h4a5f; // 0x1d44
	13'h0ea3: q2 = 16'h3c00; // 0x1d46
	13'h0ea4: q2 = 16'h4a45; // 0x1d48
	13'h0ea5: q2 = 16'h6642; // 0x1d4a
	13'h0ea6: q2 = 16'h4a79; // 0x1d4c
	13'h0ea7: q2 = 16'h0001; // 0x1d4e
	13'h0ea8: q2 = 16'h7fca; // 0x1d50
	13'h0ea9: q2 = 16'h673a; // 0x1d52
	13'h0eaa: q2 = 16'h3006; // 0x1d54
	13'h0eab: q2 = 16'h601a; // 0x1d56
	13'h0eac: q2 = 16'h4eb9; // 0x1d58
	13'h0ead: q2 = 16'h0000; // 0x1d5a
	13'h0eae: q2 = 16'ha4e4; // 0x1d5c
	13'h0eaf: q2 = 16'h6026; // 0x1d5e
	13'h0eb0: q2 = 16'h4eb9; // 0x1d60
	13'h0eb1: q2 = 16'h0000; // 0x1d62
	13'h0eb2: q2 = 16'haa5c; // 0x1d64
	13'h0eb3: q2 = 16'h601e; // 0x1d66
	13'h0eb4: q2 = 16'h4eb9; // 0x1d68
	13'h0eb5: q2 = 16'h0000; // 0x1d6a
	13'h0eb6: q2 = 16'h9da6; // 0x1d6c
	13'h0eb7: q2 = 16'h6016; // 0x1d6e
	13'h0eb8: q2 = 16'h6014; // 0x1d70
	13'h0eb9: q2 = 16'hb07c; // 0x1d72
	13'h0eba: q2 = 16'h0002; // 0x1d74
	13'h0ebb: q2 = 16'h620e; // 0x1d76
	13'h0ebc: q2 = 16'he540; // 0x1d78
	13'h0ebd: q2 = 16'h3040; // 0x1d7a
	13'h0ebe: q2 = 16'hd1fc; // 0x1d7c
	13'h0ebf: q2 = 16'h0000; // 0x1d7e
	13'h0ec0: q2 = 16'hfa06; // 0x1d80
	13'h0ec1: q2 = 16'h2050; // 0x1d82
	13'h0ec2: q2 = 16'h4ed0; // 0x1d84
	13'h0ec3: q2 = 16'h4eb9; // 0x1d86
	13'h0ec4: q2 = 16'h0000; // 0x1d88
	13'h0ec5: q2 = 16'h0226; // 0x1d8a
	13'h0ec6: q2 = 16'h7a01; // 0x1d8c
	13'h0ec7: q2 = 16'h4a79; // 0x1d8e
	13'h0ec8: q2 = 16'h0001; // 0x1d90
	13'h0ec9: q2 = 16'h7fca; // 0x1d92
	13'h0eca: q2 = 16'h6602; // 0x1d94
	13'h0ecb: q2 = 16'h4245; // 0x1d96
	13'h0ecc: q2 = 16'h6000; // 0x1d98
	13'h0ecd: q2 = 16'hff36; // 0x1d9a
	13'h0ece: q2 = 16'h4a9f; // 0x1d9c
	13'h0ecf: q2 = 16'h4cdf; // 0x1d9e
	13'h0ed0: q2 = 16'h00f8; // 0x1da0
	13'h0ed1: q2 = 16'h4e5e; // 0x1da2
	13'h0ed2: q2 = 16'h4e75; // 0x1da4
	13'h0ed3: q2 = 16'h4e56; // 0x1da6
	13'h0ed4: q2 = 16'hffd8; // 0x1da8
	13'h0ed5: q2 = 16'h48e7; // 0x1daa
	13'h0ed6: q2 = 16'h3f04; // 0x1dac
	13'h0ed7: q2 = 16'h2a7c; // 0x1dae
	13'h0ed8: q2 = 16'h0001; // 0x1db0
	13'h0ed9: q2 = 16'h86b8; // 0x1db2
	13'h0eda: q2 = 16'h4245; // 0x1db4
	13'h0edb: q2 = 16'h3d7c; // 0x1db6
	13'h0edc: q2 = 16'h0001; // 0x1db8
	13'h0edd: q2 = 16'hfffe; // 0x1dba
	13'h0ede: q2 = 16'h426e; // 0x1dbc
	13'h0edf: q2 = 16'hfffc; // 0x1dbe
	13'h0ee0: q2 = 16'h3d7c; // 0x1dc0
	13'h0ee1: q2 = 16'h0001; // 0x1dc2
	13'h0ee2: q2 = 16'hfffa; // 0x1dc4
	13'h0ee3: q2 = 16'h4eb9; // 0x1dc6
	13'h0ee4: q2 = 16'h0000; // 0x1dc8
	13'h0ee5: q2 = 16'h1564; // 0x1dca
	13'h0ee6: q2 = 16'h7e0a; // 0x1dcc
	13'h0ee7: q2 = 16'hbe7c; // 0x1dce
	13'h0ee8: q2 = 16'h000e; // 0x1dd0
	13'h0ee9: q2 = 16'h6c10; // 0x1dd2
	13'h0eea: q2 = 16'h3007; // 0x1dd4
	13'h0eeb: q2 = 16'he340; // 0x1dd6
	13'h0eec: q2 = 16'h48c0; // 0x1dd8
	13'h0eed: q2 = 16'hd08d; // 0x1dda
	13'h0eee: q2 = 16'h2040; // 0x1ddc
	13'h0eef: q2 = 16'h4250; // 0x1dde
	13'h0ef0: q2 = 16'h5247; // 0x1de0
	13'h0ef1: q2 = 16'h60ea; // 0x1de2
	13'h0ef2: q2 = 16'h4eb9; // 0x1de4
	13'h0ef3: q2 = 16'h0000; // 0x1de6
	13'h0ef4: q2 = 16'h0226; // 0x1de8
	13'h0ef5: q2 = 16'h4247; // 0x1dea
	13'h0ef6: q2 = 16'hbe7c; // 0x1dec
	13'h0ef7: q2 = 16'h0007; // 0x1dee
	13'h0ef8: q2 = 16'h6c58; // 0x1df0
	13'h0ef9: q2 = 16'hbe7c; // 0x1df2
	13'h0efa: q2 = 16'h0004; // 0x1df4
	13'h0efb: q2 = 16'h6c04; // 0x1df6
	13'h0efc: q2 = 16'h7664; // 0x1df8
	13'h0efd: q2 = 16'h6002; // 0x1dfa
	13'h0efe: q2 = 16'h4243; // 0x1dfc
	13'h0eff: q2 = 16'h3eb9; // 0x1dfe
	13'h0f00: q2 = 16'h0000; // 0x1e00
	13'h0f01: q2 = 16'hfa12; // 0x1e02
	13'h0f02: q2 = 16'h3007; // 0x1e04
	13'h0f03: q2 = 16'hd157; // 0x1e06
	13'h0f04: q2 = 16'h200e; // 0x1e08
	13'h0f05: q2 = 16'hd0bc; // 0x1e0a
	13'h0f06: q2 = 16'hffff; // 0x1e0c
	13'h0f07: q2 = 16'hffd8; // 0x1e0e
	13'h0f08: q2 = 16'h2f00; // 0x1e10
	13'h0f09: q2 = 16'h4eb9; // 0x1e12
	13'h0f0a: q2 = 16'h0000; // 0x1e14
	13'h0f0b: q2 = 16'h78f6; // 0x1e16
	13'h0f0c: q2 = 16'h4a9f; // 0x1e18
	13'h0f0d: q2 = 16'h3ebc; // 0x1e1a
	13'h0f0e: q2 = 16'h0036; // 0x1e1c
	13'h0f0f: q2 = 16'h4267; // 0x1e1e
	13'h0f10: q2 = 16'h3f03; // 0x1e20
	13'h0f11: q2 = 16'h3007; // 0x1e22
	13'h0f12: q2 = 16'he340; // 0x1e24
	13'h0f13: q2 = 16'h48c0; // 0x1e26
	13'h0f14: q2 = 16'hd0bc; // 0x1e28
	13'h0f15: q2 = 16'h0000; // 0x1e2a
	13'h0f16: q2 = 16'hfa14; // 0x1e2c
	13'h0f17: q2 = 16'h2040; // 0x1e2e
	13'h0f18: q2 = 16'h3f10; // 0x1e30
	13'h0f19: q2 = 16'h200e; // 0x1e32
	13'h0f1a: q2 = 16'hd0bc; // 0x1e34
	13'h0f1b: q2 = 16'hffff; // 0x1e36
	13'h0f1c: q2 = 16'hffd8; // 0x1e38
	13'h0f1d: q2 = 16'h2f00; // 0x1e3a
	13'h0f1e: q2 = 16'h4eb9; // 0x1e3c
	13'h0f1f: q2 = 16'h0000; // 0x1e3e
	13'h0f20: q2 = 16'h026c; // 0x1e40
	13'h0f21: q2 = 16'hdefc; // 0x1e42
	13'h0f22: q2 = 16'h000a; // 0x1e44
	13'h0f23: q2 = 16'h5247; // 0x1e46
	13'h0f24: q2 = 16'h60a2; // 0x1e48
	13'h0f25: q2 = 16'h4247; // 0x1e4a
	13'h0f26: q2 = 16'hbe7c; // 0x1e4c
	13'h0f27: q2 = 16'h000e; // 0x1e4e
	13'h0f28: q2 = 16'h6c00; // 0x1e50
	13'h0f29: q2 = 16'h016a; // 0x1e52
	13'h0f2a: q2 = 16'hbe45; // 0x1e54
	13'h0f2b: q2 = 16'h6604; // 0x1e56
	13'h0f2c: q2 = 16'h782d; // 0x1e58
	13'h0f2d: q2 = 16'h6002; // 0x1e5a
	13'h0f2e: q2 = 16'h7836; // 0x1e5c
	13'h0f2f: q2 = 16'h3eb9; // 0x1e5e
	13'h0f30: q2 = 16'h0000; // 0x1e60
	13'h0f31: q2 = 16'hfa22; // 0x1e62
	13'h0f32: q2 = 16'h3007; // 0x1e64
	13'h0f33: q2 = 16'hd157; // 0x1e66
	13'h0f34: q2 = 16'h200e; // 0x1e68
	13'h0f35: q2 = 16'hd0bc; // 0x1e6a
	13'h0f36: q2 = 16'hffff; // 0x1e6c
	13'h0f37: q2 = 16'hffd8; // 0x1e6e
	13'h0f38: q2 = 16'h2f00; // 0x1e70
	13'h0f39: q2 = 16'h4eb9; // 0x1e72
	13'h0f3a: q2 = 16'h0000; // 0x1e74
	13'h0f3b: q2 = 16'h78f6; // 0x1e76
	13'h0f3c: q2 = 16'h4a9f; // 0x1e78
	13'h0f3d: q2 = 16'h3e84; // 0x1e7a
	13'h0f3e: q2 = 16'h4267; // 0x1e7c
	13'h0f3f: q2 = 16'h3f3c; // 0x1e7e
	13'h0f40: q2 = 16'h0003; // 0x1e80
	13'h0f41: q2 = 16'h3007; // 0x1e82
	13'h0f42: q2 = 16'he340; // 0x1e84
	13'h0f43: q2 = 16'h48c0; // 0x1e86
	13'h0f44: q2 = 16'hd0bc; // 0x1e88
	13'h0f45: q2 = 16'h0000; // 0x1e8a
	13'h0f46: q2 = 16'hfa24; // 0x1e8c
	13'h0f47: q2 = 16'h2040; // 0x1e8e
	13'h0f48: q2 = 16'h3f10; // 0x1e90
	13'h0f49: q2 = 16'h200e; // 0x1e92
	13'h0f4a: q2 = 16'hd0bc; // 0x1e94
	13'h0f4b: q2 = 16'hffff; // 0x1e96
	13'h0f4c: q2 = 16'hffd8; // 0x1e98
	13'h0f4d: q2 = 16'h2f00; // 0x1e9a
	13'h0f4e: q2 = 16'h4eb9; // 0x1e9c
	13'h0f4f: q2 = 16'h0000; // 0x1e9e
	13'h0f50: q2 = 16'h026c; // 0x1ea0
	13'h0f51: q2 = 16'hdefc; // 0x1ea2
	13'h0f52: q2 = 16'h000a; // 0x1ea4
	13'h0f53: q2 = 16'hbe7c; // 0x1ea6
	13'h0f54: q2 = 16'h0009; // 0x1ea8
	13'h0f55: q2 = 16'h6f30; // 0x1eaa
	13'h0f56: q2 = 16'h3007; // 0x1eac
	13'h0f57: q2 = 16'he340; // 0x1eae
	13'h0f58: q2 = 16'h48c0; // 0x1eb0
	13'h0f59: q2 = 16'hd08d; // 0x1eb2
	13'h0f5a: q2 = 16'h2040; // 0x1eb4
	13'h0f5b: q2 = 16'h0c50; // 0x1eb6
	13'h0f5c: q2 = 16'h0002; // 0x1eb8
	13'h0f5d: q2 = 16'h6720; // 0x1eba
	13'h0f5e: q2 = 16'hbe45; // 0x1ebc
	13'h0f5f: q2 = 16'h6610; // 0x1ebe
	13'h0f60: q2 = 16'h3007; // 0x1ec0
	13'h0f61: q2 = 16'he340; // 0x1ec2
	13'h0f62: q2 = 16'h48c0; // 0x1ec4
	13'h0f63: q2 = 16'hd08d; // 0x1ec6
	13'h0f64: q2 = 16'h2040; // 0x1ec8
	13'h0f65: q2 = 16'h30bc; // 0x1eca
	13'h0f66: q2 = 16'h0001; // 0x1ecc
	13'h0f67: q2 = 16'h600c; // 0x1ece
	13'h0f68: q2 = 16'h3007; // 0x1ed0
	13'h0f69: q2 = 16'he340; // 0x1ed2
	13'h0f6a: q2 = 16'h48c0; // 0x1ed4
	13'h0f6b: q2 = 16'hd08d; // 0x1ed6
	13'h0f6c: q2 = 16'h2040; // 0x1ed8
	13'h0f6d: q2 = 16'h4250; // 0x1eda
	13'h0f6e: q2 = 16'hbe7c; // 0x1edc
	13'h0f6f: q2 = 16'h0002; // 0x1ede
	13'h0f70: q2 = 16'h6706; // 0x1ee0
	13'h0f71: q2 = 16'hbe7c; // 0x1ee2
	13'h0f72: q2 = 16'h0003; // 0x1ee4
	13'h0f73: q2 = 16'h665e; // 0x1ee6
	13'h0f74: q2 = 16'h3007; // 0x1ee8
	13'h0f75: q2 = 16'he340; // 0x1eea
	13'h0f76: q2 = 16'h48c0; // 0x1eec
	13'h0f77: q2 = 16'hd08d; // 0x1eee
	13'h0f78: q2 = 16'h2040; // 0x1ef0
	13'h0f79: q2 = 16'h3010; // 0x1ef2
	13'h0f7a: q2 = 16'hc1fc; // 0x1ef4
	13'h0f7b: q2 = 16'h0032; // 0x1ef6
	13'h0f7c: q2 = 16'h3c00; // 0x1ef8
	13'h0f7d: q2 = 16'h4a46; // 0x1efa
	13'h0f7e: q2 = 16'h672e; // 0x1efc
	13'h0f7f: q2 = 16'h200e; // 0x1efe
	13'h0f80: q2 = 16'hd0bc; // 0x1f00
	13'h0f81: q2 = 16'hffff; // 0x1f02
	13'h0f82: q2 = 16'hffd8; // 0x1f04
	13'h0f83: q2 = 16'h2e80; // 0x1f06
	13'h0f84: q2 = 16'h3f06; // 0x1f08
	13'h0f85: q2 = 16'h4eb9; // 0x1f0a
	13'h0f86: q2 = 16'h0000; // 0x1f0c
	13'h0f87: q2 = 16'h0828; // 0x1f0e
	13'h0f88: q2 = 16'h4a5f; // 0x1f10
	13'h0f89: q2 = 16'h2ebc; // 0x1f12
	13'h0f8a: q2 = 16'h0000; // 0x1f14
	13'h0f8b: q2 = 16'hfa7a; // 0x1f16
	13'h0f8c: q2 = 16'h200e; // 0x1f18
	13'h0f8d: q2 = 16'hd0bc; // 0x1f1a
	13'h0f8e: q2 = 16'hffff; // 0x1f1c
	13'h0f8f: q2 = 16'hffd8; // 0x1f1e
	13'h0f90: q2 = 16'h2f00; // 0x1f20
	13'h0f91: q2 = 16'h4eb9; // 0x1f22
	13'h0f92: q2 = 16'h0000; // 0x1f24
	13'h0f93: q2 = 16'h0770; // 0x1f26
	13'h0f94: q2 = 16'h4a9f; // 0x1f28
	13'h0f95: q2 = 16'h6018; // 0x1f2a
	13'h0f96: q2 = 16'h2ebc; // 0x1f2c
	13'h0f97: q2 = 16'h0000; // 0x1f2e
	13'h0f98: q2 = 16'hfa7d; // 0x1f30
	13'h0f99: q2 = 16'h200e; // 0x1f32
	13'h0f9a: q2 = 16'hd0bc; // 0x1f34
	13'h0f9b: q2 = 16'hffff; // 0x1f36
	13'h0f9c: q2 = 16'hffd8; // 0x1f38
	13'h0f9d: q2 = 16'h2f00; // 0x1f3a
	13'h0f9e: q2 = 16'h4eb9; // 0x1f3c
	13'h0f9f: q2 = 16'h0000; // 0x1f3e
	13'h0fa0: q2 = 16'h0750; // 0x1f40
	13'h0fa1: q2 = 16'h4a9f; // 0x1f42
	13'h0fa2: q2 = 16'h6038; // 0x1f44
	13'h0fa3: q2 = 16'h3007; // 0x1f46
	13'h0fa4: q2 = 16'he340; // 0x1f48
	13'h0fa5: q2 = 16'h48c0; // 0x1f4a
	13'h0fa6: q2 = 16'hd0bc; // 0x1f4c
	13'h0fa7: q2 = 16'h0000; // 0x1f4e
	13'h0fa8: q2 = 16'hfa5c; // 0x1f50
	13'h0fa9: q2 = 16'h2040; // 0x1f52
	13'h0faa: q2 = 16'h3e90; // 0x1f54
	13'h0fab: q2 = 16'h3007; // 0x1f56
	13'h0fac: q2 = 16'he340; // 0x1f58
	13'h0fad: q2 = 16'h48c0; // 0x1f5a
	13'h0fae: q2 = 16'hd08d; // 0x1f5c
	13'h0faf: q2 = 16'h2040; // 0x1f5e
	13'h0fb0: q2 = 16'h3010; // 0x1f60
	13'h0fb1: q2 = 16'hd157; // 0x1f62
	13'h0fb2: q2 = 16'h3039; // 0x1f64
	13'h0fb3: q2 = 16'h0000; // 0x1f66
	13'h0fb4: q2 = 16'hfa78; // 0x1f68
	13'h0fb5: q2 = 16'hd157; // 0x1f6a
	13'h0fb6: q2 = 16'h200e; // 0x1f6c
	13'h0fb7: q2 = 16'hd0bc; // 0x1f6e
	13'h0fb8: q2 = 16'hffff; // 0x1f70
	13'h0fb9: q2 = 16'hffd8; // 0x1f72
	13'h0fba: q2 = 16'h2f00; // 0x1f74
	13'h0fbb: q2 = 16'h4eb9; // 0x1f76
	13'h0fbc: q2 = 16'h0000; // 0x1f78
	13'h0fbd: q2 = 16'h78f6; // 0x1f7a
	13'h0fbe: q2 = 16'h4a9f; // 0x1f7c
	13'h0fbf: q2 = 16'hbe7c; // 0x1f7e
	13'h0fc0: q2 = 16'h0009; // 0x1f80
	13'h0fc1: q2 = 16'h6f04; // 0x1f82
	13'h0fc2: q2 = 16'h7c0a; // 0x1f84
	13'h0fc3: q2 = 16'h6002; // 0x1f86
	13'h0fc4: q2 = 16'h7c08; // 0x1f88
	13'h0fc5: q2 = 16'h3e84; // 0x1f8a
	13'h0fc6: q2 = 16'h3f06; // 0x1f8c
	13'h0fc7: q2 = 16'h3f3c; // 0x1f8e
	13'h0fc8: q2 = 16'hffe1; // 0x1f90
	13'h0fc9: q2 = 16'h3007; // 0x1f92
	13'h0fca: q2 = 16'he340; // 0x1f94
	13'h0fcb: q2 = 16'h48c0; // 0x1f96
	13'h0fcc: q2 = 16'hd0bc; // 0x1f98
	13'h0fcd: q2 = 16'h0000; // 0x1f9a
	13'h0fce: q2 = 16'hfa24; // 0x1f9c
	13'h0fcf: q2 = 16'h2040; // 0x1f9e
	13'h0fd0: q2 = 16'h3f10; // 0x1fa0
	13'h0fd1: q2 = 16'h200e; // 0x1fa2
	13'h0fd2: q2 = 16'hd0bc; // 0x1fa4
	13'h0fd3: q2 = 16'hffff; // 0x1fa6
	13'h0fd4: q2 = 16'hffd8; // 0x1fa8
	13'h0fd5: q2 = 16'h2f00; // 0x1faa
	13'h0fd6: q2 = 16'h4eb9; // 0x1fac
	13'h0fd7: q2 = 16'h0000; // 0x1fae
	13'h0fd8: q2 = 16'h026c; // 0x1fb0
	13'h0fd9: q2 = 16'hdefc; // 0x1fb2
	13'h0fda: q2 = 16'h000a; // 0x1fb4
	13'h0fdb: q2 = 16'h5247; // 0x1fb6
	13'h0fdc: q2 = 16'h6000; // 0x1fb8
	13'h0fdd: q2 = 16'hfe92; // 0x1fba
	13'h0fde: q2 = 16'h3ebc; // 0x1fbc
	13'h0fdf: q2 = 16'h000d; // 0x1fbe
	13'h0fe0: q2 = 16'h3f05; // 0x1fc0
	13'h0fe1: q2 = 16'h4eb9; // 0x1fc2
	13'h0fe2: q2 = 16'h0000; // 0x1fc4
	13'h0fe3: q2 = 16'ha602; // 0x1fc6
	13'h0fe4: q2 = 16'h4a5f; // 0x1fc8
	13'h0fe5: q2 = 16'h3a00; // 0x1fca
	13'h0fe6: q2 = 16'h4a79; // 0x1fcc
	13'h0fe7: q2 = 16'h0001; // 0x1fce
	13'h0fe8: q2 = 16'h7fca; // 0x1fd0
	13'h0fe9: q2 = 16'h6700; // 0x1fd2
	13'h0fea: q2 = 16'h0100; // 0x1fd4
	13'h0feb: q2 = 16'h4a6e; // 0x1fd6
	13'h0fec: q2 = 16'hfffa; // 0x1fd8
	13'h0fed: q2 = 16'h6600; // 0x1fda
	13'h0fee: q2 = 16'h00f8; // 0x1fdc
	13'h0fef: q2 = 16'h4ab9; // 0x1fde
	13'h0ff0: q2 = 16'h0001; // 0x1fe0
	13'h0ff1: q2 = 16'h7fc2; // 0x1fe2
	13'h0ff2: q2 = 16'h6f08; // 0x1fe4
	13'h0ff3: q2 = 16'h4a6e; // 0x1fe6
	13'h0ff4: q2 = 16'hfffc; // 0x1fe8
	13'h0ff5: q2 = 16'h6600; // 0x1fea
	13'h0ff6: q2 = 16'h00e8; // 0x1fec
	13'h0ff7: q2 = 16'hba7c; // 0x1fee
	13'h0ff8: q2 = 16'h000a; // 0x1ff0
	13'h0ff9: q2 = 16'h6c00; // 0x1ff2
	13'h0ffa: q2 = 16'h008a; // 0x1ff4
	13'h0ffb: q2 = 16'h3005; // 0x1ff6
	13'h0ffc: q2 = 16'he340; // 0x1ff8
	13'h0ffd: q2 = 16'h48c0; // 0x1ffa
	13'h0ffe: q2 = 16'hd08d; // 0x1ffc
	13'h0fff: q2 = 16'h2040; // 0x1ffe
	13'h1000: q2 = 16'h5250; // 0x2000
	13'h1001: q2 = 16'h3005; // 0x2002
	13'h1002: q2 = 16'he340; // 0x2004
	13'h1003: q2 = 16'h48c0; // 0x2006
	13'h1004: q2 = 16'hd08d; // 0x2008
	13'h1005: q2 = 16'h2040; // 0x200a
	13'h1006: q2 = 16'h3010; // 0x200c
	13'h1007: q2 = 16'h3205; // 0x200e
	13'h1008: q2 = 16'he341; // 0x2010
	13'h1009: q2 = 16'h48c1; // 0x2012
	13'h100a: q2 = 16'hd2bc; // 0x2014
	13'h100b: q2 = 16'h0000; // 0x2016
	13'h100c: q2 = 16'hfa40; // 0x2018
	13'h100d: q2 = 16'h2241; // 0x201a
	13'h100e: q2 = 16'hb051; // 0x201c
	13'h100f: q2 = 16'h6d0c; // 0x201e
	13'h1010: q2 = 16'h3005; // 0x2020
	13'h1011: q2 = 16'he340; // 0x2022
	13'h1012: q2 = 16'h48c0; // 0x2024
	13'h1013: q2 = 16'hd08d; // 0x2026
	13'h1014: q2 = 16'h2040; // 0x2028
	13'h1015: q2 = 16'h4250; // 0x202a
	13'h1016: q2 = 16'hba7c; // 0x202c
	13'h1017: q2 = 16'h0002; // 0x202e
	13'h1018: q2 = 16'h661c; // 0x2030
	13'h1019: q2 = 16'h4a79; // 0x2032
	13'h101a: q2 = 16'h0001; // 0x2034
	13'h101b: q2 = 16'h86be; // 0x2036
	13'h101c: q2 = 16'h6714; // 0x2038
	13'h101d: q2 = 16'h3039; // 0x203a
	13'h101e: q2 = 16'h0001; // 0x203c
	13'h101f: q2 = 16'h86bc; // 0x203e
	13'h1020: q2 = 16'hb079; // 0x2040
	13'h1021: q2 = 16'h0001; // 0x2042
	13'h1022: q2 = 16'h86be; // 0x2044
	13'h1023: q2 = 16'h6f06; // 0x2046
	13'h1024: q2 = 16'h4279; // 0x2048
	13'h1025: q2 = 16'h0001; // 0x204a
	13'h1026: q2 = 16'h86bc; // 0x204c
	13'h1027: q2 = 16'hba7c; // 0x204e
	13'h1028: q2 = 16'h0003; // 0x2050
	13'h1029: q2 = 16'h661c; // 0x2052
	13'h102a: q2 = 16'h4a79; // 0x2054
	13'h102b: q2 = 16'h0001; // 0x2056
	13'h102c: q2 = 16'h86bc; // 0x2058
	13'h102d: q2 = 16'h6714; // 0x205a
	13'h102e: q2 = 16'h0c79; // 0x205c
	13'h102f: q2 = 16'h0001; // 0x205e
	13'h1030: q2 = 16'h0001; // 0x2060
	13'h1031: q2 = 16'h86be; // 0x2062
	13'h1032: q2 = 16'h660a; // 0x2064
	13'h1033: q2 = 16'h33f9; // 0x2066
	13'h1034: q2 = 16'h0001; // 0x2068
	13'h1035: q2 = 16'h86bc; // 0x206a
	13'h1036: q2 = 16'h0001; // 0x206c
	13'h1037: q2 = 16'h86be; // 0x206e
	13'h1038: q2 = 16'h4279; // 0x2070
	13'h1039: q2 = 16'h0001; // 0x2072
	13'h103a: q2 = 16'h86cc; // 0x2074
	13'h103b: q2 = 16'h4279; // 0x2076
	13'h103c: q2 = 16'h0001; // 0x2078
	13'h103d: q2 = 16'h86ce; // 0x207a
	13'h103e: q2 = 16'h600e; // 0x207c
	13'h103f: q2 = 16'h3005; // 0x207e
	13'h1040: q2 = 16'he340; // 0x2080
	13'h1041: q2 = 16'h48c0; // 0x2082
	13'h1042: q2 = 16'hd08d; // 0x2084
	13'h1043: q2 = 16'h2040; // 0x2086
	13'h1044: q2 = 16'h30bc; // 0x2088
	13'h1045: q2 = 16'h0002; // 0x208a
	13'h1046: q2 = 16'hba7c; // 0x208c
	13'h1047: q2 = 16'h000a; // 0x208e
	13'h1048: q2 = 16'h660c; // 0x2090
	13'h1049: q2 = 16'h4eb9; // 0x2092
	13'h104a: q2 = 16'h0000; // 0x2094
	13'h104b: q2 = 16'h1564; // 0x2096
	13'h104c: q2 = 16'h4279; // 0x2098
	13'h104d: q2 = 16'h0001; // 0x209a
	13'h104e: q2 = 16'h86ce; // 0x209c
	13'h104f: q2 = 16'hba7c; // 0x209e
	13'h1050: q2 = 16'h000b; // 0x20a0
	13'h1051: q2 = 16'h660c; // 0x20a2
	13'h1052: q2 = 16'h4eb9; // 0x20a4
	13'h1053: q2 = 16'h0000; // 0x20a6
	13'h1054: q2 = 16'h3cda; // 0x20a8
	13'h1055: q2 = 16'h4279; // 0x20aa
	13'h1056: q2 = 16'h0001; // 0x20ac
	13'h1057: q2 = 16'h86cc; // 0x20ae
	13'h1058: q2 = 16'h4a6e; // 0x20b0
	13'h1059: q2 = 16'hfffc; // 0x20b2
	13'h105a: q2 = 16'h670c; // 0x20b4
	13'h105b: q2 = 16'h23fc; // 0x20b6
	13'h105c: q2 = 16'h0000; // 0x20b8
	13'h105d: q2 = 16'h0004; // 0x20ba
	13'h105e: q2 = 16'h0001; // 0x20bc
	13'h105f: q2 = 16'h7fc2; // 0x20be
	13'h1060: q2 = 16'h6010; // 0x20c0
	13'h1061: q2 = 16'h23fc; // 0x20c2
	13'h1062: q2 = 16'h0000; // 0x20c4
	13'h1063: q2 = 16'h0028; // 0x20c6
	13'h1064: q2 = 16'h0001; // 0x20c8
	13'h1065: q2 = 16'h7fc2; // 0x20ca
	13'h1066: q2 = 16'h3d7c; // 0x20cc
	13'h1067: q2 = 16'h0001; // 0x20ce
	13'h1068: q2 = 16'hfffc; // 0x20d0
	13'h1069: q2 = 16'h6010; // 0x20d2
	13'h106a: q2 = 16'h4a79; // 0x20d4
	13'h106b: q2 = 16'h0001; // 0x20d6
	13'h106c: q2 = 16'h7fca; // 0x20d8
	13'h106d: q2 = 16'h6608; // 0x20da
	13'h106e: q2 = 16'h426e; // 0x20dc
	13'h106f: q2 = 16'hfffc; // 0x20de
	13'h1070: q2 = 16'h426e; // 0x20e0
	13'h1071: q2 = 16'hfffa; // 0x20e2
	13'h1072: q2 = 16'h4a79; // 0x20e4
	13'h1073: q2 = 16'h0001; // 0x20e6
	13'h1074: q2 = 16'h8a7e; // 0x20e8
	13'h1075: q2 = 16'h6604; // 0x20ea
	13'h1076: q2 = 16'h426e; // 0x20ec
	13'h1077: q2 = 16'hfffe; // 0x20ee
	13'h1078: q2 = 16'h4a6e; // 0x20f0
	13'h1079: q2 = 16'hfffe; // 0x20f2
	13'h107a: q2 = 16'h6632; // 0x20f4
	13'h107b: q2 = 16'h4a79; // 0x20f6
	13'h107c: q2 = 16'h0001; // 0x20f8
	13'h107d: q2 = 16'h8a7e; // 0x20fa
	13'h107e: q2 = 16'h672a; // 0x20fc
	13'h107f: q2 = 16'h4eb9; // 0x20fe
	13'h1080: q2 = 16'h0000; // 0x2100
	13'h1081: q2 = 16'hb2ae; // 0x2102
	13'h1082: q2 = 16'h0c79; // 0x2104
	13'h1083: q2 = 16'h0002; // 0x2106
	13'h1084: q2 = 16'h0001; // 0x2108
	13'h1085: q2 = 16'h86d0; // 0x210a
	13'h1086: q2 = 16'h6608; // 0x210c
	13'h1087: q2 = 16'h4257; // 0x210e
	13'h1088: q2 = 16'h4eb9; // 0x2110
	13'h1089: q2 = 16'h0000; // 0x2112
	13'h108a: q2 = 16'h55ce; // 0x2114
	13'h108b: q2 = 16'h0c79; // 0x2116
	13'h108c: q2 = 16'h0002; // 0x2118
	13'h108d: q2 = 16'h0001; // 0x211a
	13'h108e: q2 = 16'h86d2; // 0x211c
	13'h108f: q2 = 16'h6606; // 0x211e
	13'h1090: q2 = 16'h4eb9; // 0x2120
	13'h1091: q2 = 16'h0000; // 0x2122
	13'h1092: q2 = 16'haa34; // 0x2124
	13'h1093: q2 = 16'h6004; // 0x2126
	13'h1094: q2 = 16'h6000; // 0x2128
	13'h1095: q2 = 16'hfd20; // 0x212a
	13'h1096: q2 = 16'h4a9f; // 0x212c
	13'h1097: q2 = 16'h4cdf; // 0x212e
	13'h1098: q2 = 16'h20f8; // 0x2130
	13'h1099: q2 = 16'h4e5e; // 0x2132
	13'h109a: q2 = 16'h4e75; // 0x2134
	13'h109b: q2 = 16'h4e56; // 0x2136
	13'h109c: q2 = 16'hffde; // 0x2138
	13'h109d: q2 = 16'h48e7; // 0x213a
	13'h109e: q2 = 16'h0700; // 0x213c
	13'h109f: q2 = 16'h4eb9; // 0x213e
	13'h10a0: q2 = 16'h0000; // 0x2140
	13'h10a1: q2 = 16'h0226; // 0x2142
	13'h10a2: q2 = 16'h4247; // 0x2144
	13'h10a3: q2 = 16'hbe7c; // 0x2146
	13'h10a4: q2 = 16'h0002; // 0x2148
	13'h10a5: q2 = 16'h6e4e; // 0x214a
	13'h10a6: q2 = 16'h3eb9; // 0x214c
	13'h10a7: q2 = 16'h0000; // 0x214e
	13'h10a8: q2 = 16'hf9dc; // 0x2150
	13'h10a9: q2 = 16'h3007; // 0x2152
	13'h10aa: q2 = 16'hd157; // 0x2154
	13'h10ab: q2 = 16'h200e; // 0x2156
	13'h10ac: q2 = 16'hd0bc; // 0x2158
	13'h10ad: q2 = 16'hffff; // 0x215a
	13'h10ae: q2 = 16'hffde; // 0x215c
	13'h10af: q2 = 16'h2f00; // 0x215e
	13'h10b0: q2 = 16'h4eb9; // 0x2160
	13'h10b1: q2 = 16'h0000; // 0x2162
	13'h10b2: q2 = 16'h78f6; // 0x2164
	13'h10b3: q2 = 16'h4a9f; // 0x2166
	13'h10b4: q2 = 16'h3ebc; // 0x2168
	13'h10b5: q2 = 16'h0036; // 0x216a
	13'h10b6: q2 = 16'h4267; // 0x216c
	13'h10b7: q2 = 16'h3f3c; // 0x216e
	13'h10b8: q2 = 16'h0064; // 0x2170
	13'h10b9: q2 = 16'h3007; // 0x2172
	13'h10ba: q2 = 16'he340; // 0x2174
	13'h10bb: q2 = 16'h48c0; // 0x2176
	13'h10bc: q2 = 16'hd0bc; // 0x2178
	13'h10bd: q2 = 16'h0000; // 0x217a
	13'h10be: q2 = 16'hf9de; // 0x217c
	13'h10bf: q2 = 16'h2040; // 0x217e
	13'h10c0: q2 = 16'h3f10; // 0x2180
	13'h10c1: q2 = 16'h200e; // 0x2182
	13'h10c2: q2 = 16'hd0bc; // 0x2184
	13'h10c3: q2 = 16'hffff; // 0x2186
	13'h10c4: q2 = 16'hffde; // 0x2188
	13'h10c5: q2 = 16'h2f00; // 0x218a
	13'h10c6: q2 = 16'h4eb9; // 0x218c
	13'h10c7: q2 = 16'h0000; // 0x218e
	13'h10c8: q2 = 16'h026c; // 0x2190
	13'h10c9: q2 = 16'hdefc; // 0x2192
	13'h10ca: q2 = 16'h000a; // 0x2194
	13'h10cb: q2 = 16'h5247; // 0x2196
	13'h10cc: q2 = 16'h60ac; // 0x2198
	13'h10cd: q2 = 16'h7c01; // 0x219a
	13'h10ce: q2 = 16'h7e01; // 0x219c
	13'h10cf: q2 = 16'h200e; // 0x219e
	13'h10d0: q2 = 16'hd0bc; // 0x21a0
	13'h10d1: q2 = 16'hffff; // 0x21a2
	13'h10d2: q2 = 16'hffde; // 0x21a4
	13'h10d3: q2 = 16'h2e80; // 0x21a6
	13'h10d4: q2 = 16'h3f07; // 0x21a8
	13'h10d5: q2 = 16'h4eb9; // 0x21aa
	13'h10d6: q2 = 16'h0000; // 0x21ac
	13'h10d7: q2 = 16'h0828; // 0x21ae
	13'h10d8: q2 = 16'h4a5f; // 0x21b0
	13'h10d9: q2 = 16'h3ebc; // 0x21b2
	13'h10da: q2 = 16'h0036; // 0x21b4
	13'h10db: q2 = 16'h3f3c; // 0x21b6
	13'h10dc: q2 = 16'h0002; // 0x21b8
	13'h10dd: q2 = 16'h3f3c; // 0x21ba
	13'h10de: q2 = 16'hffec; // 0x21bc
	13'h10df: q2 = 16'h3f3c; // 0x21be
	13'h10e0: q2 = 16'h0014; // 0x21c0
	13'h10e1: q2 = 16'h200e; // 0x21c2
	13'h10e2: q2 = 16'hd0bc; // 0x21c4
	13'h10e3: q2 = 16'hffff; // 0x21c6
	13'h10e4: q2 = 16'hffde; // 0x21c8
	13'h10e5: q2 = 16'h2f00; // 0x21ca
	13'h10e6: q2 = 16'h4eb9; // 0x21cc
	13'h10e7: q2 = 16'h0000; // 0x21ce
	13'h10e8: q2 = 16'h026c; // 0x21d0
	13'h10e9: q2 = 16'hdefc; // 0x21d2
	13'h10ea: q2 = 16'h000a; // 0x21d4
	13'h10eb: q2 = 16'h2ebc; // 0x21d6
	13'h10ec: q2 = 16'h0000; // 0x21d8
	13'h10ed: q2 = 16'hfd92; // 0x21da
	13'h10ee: q2 = 16'h4eb9; // 0x21dc
	13'h10ef: q2 = 16'h0000; // 0x21de
	13'h10f0: q2 = 16'h7e06; // 0x21e0
	13'h10f1: q2 = 16'h23fc; // 0x21e2
	13'h10f2: q2 = 16'h0000; // 0x21e4
	13'h10f3: q2 = 16'h003c; // 0x21e6
	13'h10f4: q2 = 16'h0001; // 0x21e8
	13'h10f5: q2 = 16'h7fc2; // 0x21ea
	13'h10f6: q2 = 16'h4ab9; // 0x21ec
	13'h10f7: q2 = 16'h0001; // 0x21ee
	13'h10f8: q2 = 16'h7fc2; // 0x21f0
	13'h10f9: q2 = 16'h6718; // 0x21f2
	13'h10fa: q2 = 16'h4a46; // 0x21f4
	13'h10fb: q2 = 16'h6608; // 0x21f6
	13'h10fc: q2 = 16'h4a79; // 0x21f8
	13'h10fd: q2 = 16'h0001; // 0x21fa
	13'h10fe: q2 = 16'h8a7e; // 0x21fc
	13'h10ff: q2 = 16'h660c; // 0x21fe
	13'h1100: q2 = 16'h4a79; // 0x2200
	13'h1101: q2 = 16'h0001; // 0x2202
	13'h1102: q2 = 16'h8a7e; // 0x2204
	13'h1103: q2 = 16'h6602; // 0x2206
	13'h1104: q2 = 16'h4246; // 0x2208
	13'h1105: q2 = 16'h60e0; // 0x220a
	13'h1106: q2 = 16'h4a46; // 0x220c
	13'h1107: q2 = 16'h6608; // 0x220e
	13'h1108: q2 = 16'h4a79; // 0x2210
	13'h1109: q2 = 16'h0001; // 0x2212
	13'h110a: q2 = 16'h8a7e; // 0x2214
	13'h110b: q2 = 16'h6622; // 0x2216
	13'h110c: q2 = 16'h5247; // 0x2218
	13'h110d: q2 = 16'hbe7c; // 0x221a
	13'h110e: q2 = 16'h000c; // 0x221c
	13'h110f: q2 = 16'h6f16; // 0x221e
	13'h1110: q2 = 16'h7e01; // 0x2220
	13'h1111: q2 = 16'h4279; // 0x2222
	13'h1112: q2 = 16'h0001; // 0x2224
	13'h1113: q2 = 16'h8a7a; // 0x2226
	13'h1114: q2 = 16'h4eb9; // 0x2228
	13'h1115: q2 = 16'h0000; // 0x222a
	13'h1116: q2 = 16'h8902; // 0x222c
	13'h1117: q2 = 16'h33fc; // 0x222e
	13'h1118: q2 = 16'h0001; // 0x2230
	13'h1119: q2 = 16'h0001; // 0x2232
	13'h111a: q2 = 16'h8a7a; // 0x2234
	13'h111b: q2 = 16'h6000; // 0x2236
	13'h111c: q2 = 16'hff66; // 0x2238
	13'h111d: q2 = 16'h4279; // 0x223a
	13'h111e: q2 = 16'h0001; // 0x223c
	13'h111f: q2 = 16'h8a7a; // 0x223e
	13'h1120: q2 = 16'h4eb9; // 0x2240
	13'h1121: q2 = 16'h0000; // 0x2242
	13'h1122: q2 = 16'h8902; // 0x2244
	13'h1123: q2 = 16'h33fc; // 0x2246
	13'h1124: q2 = 16'h0001; // 0x2248
	13'h1125: q2 = 16'h0001; // 0x224a
	13'h1126: q2 = 16'h8a7a; // 0x224c
	13'h1127: q2 = 16'h4a9f; // 0x224e
	13'h1128: q2 = 16'h4cdf; // 0x2250
	13'h1129: q2 = 16'h00c0; // 0x2252
	13'h112a: q2 = 16'h4e5e; // 0x2254
	13'h112b: q2 = 16'h4e75; // 0x2256
	13'h112c: q2 = 16'h4e56; // 0x2258
	13'h112d: q2 = 16'hffd8; // 0x225a
	13'h112e: q2 = 16'h48e7; // 0x225c
	13'h112f: q2 = 16'h3f0c; // 0x225e
	13'h1130: q2 = 16'h2d79; // 0x2260
	13'h1131: q2 = 16'h0000; // 0x2262
	13'h1132: q2 = 16'hfa82; // 0x2264
	13'h1133: q2 = 16'hfffa; // 0x2266
	13'h1134: q2 = 16'h4eb9; // 0x2268
	13'h1135: q2 = 16'h0000; // 0x226a
	13'h1136: q2 = 16'h0226; // 0x226c
	13'h1137: q2 = 16'h4247; // 0x226e
	13'h1138: q2 = 16'hbe7c; // 0x2270
	13'h1139: q2 = 16'h000f; // 0x2272
	13'h113a: q2 = 16'h6e6a; // 0x2274
	13'h113b: q2 = 16'hbe7c; // 0x2276
	13'h113c: q2 = 16'h0001; // 0x2278
	13'h113d: q2 = 16'h6e04; // 0x227a
	13'h113e: q2 = 16'h7c64; // 0x227c
	13'h113f: q2 = 16'h6014; // 0x227e
	13'h1140: q2 = 16'hbe7c; // 0x2280
	13'h1141: q2 = 16'h000c; // 0x2282
	13'h1142: q2 = 16'h6d0c; // 0x2284
	13'h1143: q2 = 16'h4a79; // 0x2286
	13'h1144: q2 = 16'h0001; // 0x2288
	13'h1145: q2 = 16'h758e; // 0x228a
	13'h1146: q2 = 16'h674e; // 0x228c
	13'h1147: q2 = 16'h7c10; // 0x228e
	13'h1148: q2 = 16'h6002; // 0x2290
	13'h1149: q2 = 16'h4246; // 0x2292
	13'h114a: q2 = 16'h3eb9; // 0x2294
	13'h114b: q2 = 16'h0000; // 0x2296
	13'h114c: q2 = 16'hf9e4; // 0x2298
	13'h114d: q2 = 16'h3007; // 0x229a
	13'h114e: q2 = 16'hd157; // 0x229c
	13'h114f: q2 = 16'h200e; // 0x229e
	13'h1150: q2 = 16'hd0bc; // 0x22a0
	13'h1151: q2 = 16'hffff; // 0x22a2
	13'h1152: q2 = 16'hffd8; // 0x22a4
	13'h1153: q2 = 16'h2f00; // 0x22a6
	13'h1154: q2 = 16'h4eb9; // 0x22a8
	13'h1155: q2 = 16'h0000; // 0x22aa
	13'h1156: q2 = 16'h78f6; // 0x22ac
	13'h1157: q2 = 16'h4a9f; // 0x22ae
	13'h1158: q2 = 16'h3ebc; // 0x22b0
	13'h1159: q2 = 16'h0036; // 0x22b2
	13'h115a: q2 = 16'h4267; // 0x22b4
	13'h115b: q2 = 16'h3f06; // 0x22b6
	13'h115c: q2 = 16'h3007; // 0x22b8
	13'h115d: q2 = 16'he340; // 0x22ba
	13'h115e: q2 = 16'h48c0; // 0x22bc
	13'h115f: q2 = 16'hd0bc; // 0x22be
	13'h1160: q2 = 16'h0000; // 0x22c0
	13'h1161: q2 = 16'hf9e6; // 0x22c2
	13'h1162: q2 = 16'h2040; // 0x22c4
	13'h1163: q2 = 16'h3f10; // 0x22c6
	13'h1164: q2 = 16'h200e; // 0x22c8
	13'h1165: q2 = 16'hd0bc; // 0x22ca
	13'h1166: q2 = 16'hffff; // 0x22cc
	13'h1167: q2 = 16'hffd8; // 0x22ce
	13'h1168: q2 = 16'h2f00; // 0x22d0
	13'h1169: q2 = 16'h4eb9; // 0x22d2
	13'h116a: q2 = 16'h0000; // 0x22d4
	13'h116b: q2 = 16'h026c; // 0x22d6
	13'h116c: q2 = 16'hdefc; // 0x22d8
	13'h116d: q2 = 16'h000a; // 0x22da
	13'h116e: q2 = 16'h5247; // 0x22dc
	13'h116f: q2 = 16'h6090; // 0x22de
	13'h1170: q2 = 16'h426e; // 0x22e0
	13'h1171: q2 = 16'hfffe; // 0x22e2
	13'h1172: q2 = 16'h2a7c; // 0x22e4
	13'h1173: q2 = 16'h0001; // 0x22e6
	13'h1174: q2 = 16'h8052; // 0x22e8
	13'h1175: q2 = 16'h4255; // 0x22ea
	13'h1176: q2 = 16'h287c; // 0x22ec
	13'h1177: q2 = 16'h0001; // 0x22ee
	13'h1178: q2 = 16'h7fcc; // 0x22f0
	13'h1179: q2 = 16'h206e; // 0x22f2
	13'h117a: q2 = 16'hfffa; // 0x22f4
	13'h117b: q2 = 16'h3a10; // 0x22f6
	13'h117c: q2 = 16'h7e02; // 0x22f8
	13'h117d: q2 = 16'hbe7c; // 0x22fa
	13'h117e: q2 = 16'h000f; // 0x22fc
	13'h117f: q2 = 16'h6e00; // 0x22fe
	13'h1180: q2 = 16'h01a4; // 0x2300
	13'h1181: q2 = 16'hbe7c; // 0x2302
	13'h1182: q2 = 16'h0005; // 0x2304
	13'h1183: q2 = 16'h6700; // 0x2306
	13'h1184: q2 = 16'h0196; // 0x2308
	13'h1185: q2 = 16'hbe7c; // 0x230a
	13'h1186: q2 = 16'h000d; // 0x230c
	13'h1187: q2 = 16'h6700; // 0x230e
	13'h1188: q2 = 16'h018e; // 0x2310
	13'h1189: q2 = 16'h4a79; // 0x2312
	13'h118a: q2 = 16'h0001; // 0x2314
	13'h118b: q2 = 16'h758e; // 0x2316
	13'h118c: q2 = 16'h6608; // 0x2318
	13'h118d: q2 = 16'hbe7c; // 0x231a
	13'h118e: q2 = 16'h000c; // 0x231c
	13'h118f: q2 = 16'h6c00; // 0x231e
	13'h1190: q2 = 16'h017e; // 0x2320
	13'h1191: q2 = 16'h3007; // 0x2322
	13'h1192: q2 = 16'h6000; // 0x2324
	13'h1193: q2 = 16'h00a0; // 0x2326
	13'h1194: q2 = 16'h0805; // 0x2328
	13'h1195: q2 = 16'h0002; // 0x232a
	13'h1196: q2 = 16'h6704; // 0x232c
	13'h1197: q2 = 16'h4240; // 0x232e
	13'h1198: q2 = 16'h6002; // 0x2330
	13'h1199: q2 = 16'h7001; // 0x2332
	13'h119a: q2 = 16'h3c00; // 0x2334
	13'h119b: q2 = 16'h6000; // 0x2336
	13'h119c: q2 = 16'h00a4; // 0x2338
	13'h119d: q2 = 16'h0805; // 0x233a
	13'h119e: q2 = 16'h0003; // 0x233c
	13'h119f: q2 = 16'h6704; // 0x233e
	13'h11a0: q2 = 16'h4240; // 0x2340
	13'h11a1: q2 = 16'h6002; // 0x2342
	13'h11a2: q2 = 16'h7001; // 0x2344
	13'h11a3: q2 = 16'h3c00; // 0x2346
	13'h11a4: q2 = 16'h6000; // 0x2348
	13'h11a5: q2 = 16'h0092; // 0x234a
	13'h11a6: q2 = 16'h0805; // 0x234c
	13'h11a7: q2 = 16'h0005; // 0x234e
	13'h11a8: q2 = 16'h6704; // 0x2350
	13'h11a9: q2 = 16'h4240; // 0x2352
	13'h11aa: q2 = 16'h6002; // 0x2354
	13'h11ab: q2 = 16'h7001; // 0x2356
	13'h11ac: q2 = 16'h3c00; // 0x2358
	13'h11ad: q2 = 16'h6000; // 0x235a
	13'h11ae: q2 = 16'h0080; // 0x235c
	13'h11af: q2 = 16'h3c39; // 0x235e
	13'h11b0: q2 = 16'h0001; // 0x2360
	13'h11b1: q2 = 16'h86b2; // 0x2362
	13'h11b2: q2 = 16'h6000; // 0x2364
	13'h11b3: q2 = 16'h0076; // 0x2366
	13'h11b4: q2 = 16'h3c39; // 0x2368
	13'h11b5: q2 = 16'h0001; // 0x236a
	13'h11b6: q2 = 16'h86b6; // 0x236c
	13'h11b7: q2 = 16'h6000; // 0x236e
	13'h11b8: q2 = 16'h006c; // 0x2370
	13'h11b9: q2 = 16'h0805; // 0x2372
	13'h11ba: q2 = 16'h0000; // 0x2374
	13'h11bb: q2 = 16'h6704; // 0x2376
	13'h11bc: q2 = 16'h4240; // 0x2378
	13'h11bd: q2 = 16'h6002; // 0x237a
	13'h11be: q2 = 16'h7001; // 0x237c
	13'h11bf: q2 = 16'h3c00; // 0x237e
	13'h11c0: q2 = 16'h605a; // 0x2380
	13'h11c1: q2 = 16'h0805; // 0x2382
	13'h11c2: q2 = 16'h0001; // 0x2384
	13'h11c3: q2 = 16'h6704; // 0x2386
	13'h11c4: q2 = 16'h4240; // 0x2388
	13'h11c5: q2 = 16'h6002; // 0x238a
	13'h11c6: q2 = 16'h7001; // 0x238c
	13'h11c7: q2 = 16'h3c00; // 0x238e
	13'h11c8: q2 = 16'h604a; // 0x2390
	13'h11c9: q2 = 16'h0805; // 0x2392
	13'h11ca: q2 = 16'h0004; // 0x2394
	13'h11cb: q2 = 16'h6704; // 0x2396
	13'h11cc: q2 = 16'h4240; // 0x2398
	13'h11cd: q2 = 16'h6002; // 0x239a
	13'h11ce: q2 = 16'h7001; // 0x239c
	13'h11cf: q2 = 16'h3c00; // 0x239e
	13'h11d0: q2 = 16'h603a; // 0x23a0
	13'h11d1: q2 = 16'h6038; // 0x23a2
	13'h11d2: q2 = 16'h0805; // 0x23a4
	13'h11d3: q2 = 16'h0006; // 0x23a6
	13'h11d4: q2 = 16'h6704; // 0x23a8
	13'h11d5: q2 = 16'h4240; // 0x23aa
	13'h11d6: q2 = 16'h6002; // 0x23ac
	13'h11d7: q2 = 16'h7001; // 0x23ae
	13'h11d8: q2 = 16'h3c00; // 0x23b0
	13'h11d9: q2 = 16'h6028; // 0x23b2
	13'h11da: q2 = 16'h3c39; // 0x23b4
	13'h11db: q2 = 16'h0001; // 0x23b6
	13'h11dc: q2 = 16'h86b4; // 0x23b8
	13'h11dd: q2 = 16'h6020; // 0x23ba
	13'h11de: q2 = 16'h3c39; // 0x23bc
	13'h11df: q2 = 16'h0001; // 0x23be
	13'h11e0: q2 = 16'h86da; // 0x23c0
	13'h11e1: q2 = 16'h6018; // 0x23c2
	13'h11e2: q2 = 16'h6016; // 0x23c4
	13'h11e3: q2 = 16'h5540; // 0x23c6
	13'h11e4: q2 = 16'hb07c; // 0x23c8
	13'h11e5: q2 = 16'h000d; // 0x23ca
	13'h11e6: q2 = 16'h620e; // 0x23cc
	13'h11e7: q2 = 16'he540; // 0x23ce
	13'h11e8: q2 = 16'h3040; // 0x23d0
	13'h11e9: q2 = 16'hd1fc; // 0x23d2
	13'h11ea: q2 = 16'h0000; // 0x23d4
	13'h11eb: q2 = 16'hfa86; // 0x23d6
	13'h11ec: q2 = 16'h2050; // 0x23d8
	13'h11ed: q2 = 16'h4ed0; // 0x23da
	13'h11ee: q2 = 16'hbe7c; // 0x23dc
	13'h11ef: q2 = 16'h000b; // 0x23de
	13'h11f0: q2 = 16'h6d04; // 0x23e0
	13'h11f1: q2 = 16'h761d; // 0x23e2
	13'h11f2: q2 = 16'h6002; // 0x23e4
	13'h11f3: q2 = 16'h760d; // 0x23e6
	13'h11f4: q2 = 16'hbe7c; // 0x23e8
	13'h11f5: q2 = 16'h0006; // 0x23ea
	13'h11f6: q2 = 16'h6712; // 0x23ec
	13'h11f7: q2 = 16'hbe7c; // 0x23ee
	13'h11f8: q2 = 16'h0007; // 0x23f0
	13'h11f9: q2 = 16'h670c; // 0x23f2
	13'h11fa: q2 = 16'hbe7c; // 0x23f4
	13'h11fb: q2 = 16'h000e; // 0x23f6
	13'h11fc: q2 = 16'h6706; // 0x23f8
	13'h11fd: q2 = 16'hbe7c; // 0x23fa
	13'h11fe: q2 = 16'h000f; // 0x23fc
	13'h11ff: q2 = 16'h663a; // 0x23fe
	13'h1200: q2 = 16'h4244; // 0x2400
	13'h1201: q2 = 16'hb87c; // 0x2402
	13'h1202: q2 = 16'h0008; // 0x2404
	13'h1203: q2 = 16'h6c30; // 0x2406
	13'h1204: q2 = 16'h3ebc; // 0x2408
	13'h1205: q2 = 16'h003e; // 0x240a
	13'h1206: q2 = 16'h3f06; // 0x240c
	13'h1207: q2 = 16'h0257; // 0x240e
	13'h1208: q2 = 16'h0001; // 0x2410
	13'h1209: q2 = 16'h0657; // 0x2412
	13'h120a: q2 = 16'h0030; // 0x2414
	13'h120b: q2 = 16'h3007; // 0x2416
	13'h120c: q2 = 16'he340; // 0x2418
	13'h120d: q2 = 16'h48c0; // 0x241a
	13'h120e: q2 = 16'hd0bc; // 0x241c
	13'h120f: q2 = 16'h0000; // 0x241e
	13'h1210: q2 = 16'hf9e6; // 0x2420
	13'h1211: q2 = 16'h2040; // 0x2422
	13'h1212: q2 = 16'h3f10; // 0x2424
	13'h1213: q2 = 16'h3f03; // 0x2426
	13'h1214: q2 = 16'h4eb9; // 0x2428
	13'h1215: q2 = 16'h0000; // 0x242a
	13'h1216: q2 = 16'h3d18; // 0x242c
	13'h1217: q2 = 16'h5c4f; // 0x242e
	13'h1218: q2 = 16'he246; // 0x2430
	13'h1219: q2 = 16'h5343; // 0x2432
	13'h121a: q2 = 16'h5244; // 0x2434
	13'h121b: q2 = 16'h60ca; // 0x2436
	13'h121c: q2 = 16'h6064; // 0x2438
	13'h121d: q2 = 16'hbe7c; // 0x243a
	13'h121e: q2 = 16'h000b; // 0x243c
	13'h121f: q2 = 16'h672c; // 0x243e
	13'h1220: q2 = 16'h4a46; // 0x2440
	13'h1221: q2 = 16'h6702; // 0x2442
	13'h1222: q2 = 16'h7c01; // 0x2444
	13'h1223: q2 = 16'h3ebc; // 0x2446
	13'h1224: q2 = 16'h003e; // 0x2448
	13'h1225: q2 = 16'h3f06; // 0x244a
	13'h1226: q2 = 16'h0657; // 0x244c
	13'h1227: q2 = 16'h0030; // 0x244e
	13'h1228: q2 = 16'h3007; // 0x2450
	13'h1229: q2 = 16'he340; // 0x2452
	13'h122a: q2 = 16'h48c0; // 0x2454
	13'h122b: q2 = 16'hd0bc; // 0x2456
	13'h122c: q2 = 16'h0000; // 0x2458
	13'h122d: q2 = 16'hf9e6; // 0x245a
	13'h122e: q2 = 16'h2040; // 0x245c
	13'h122f: q2 = 16'h3f10; // 0x245e
	13'h1230: q2 = 16'h3f03; // 0x2460
	13'h1231: q2 = 16'h4eb9; // 0x2462
	13'h1232: q2 = 16'h0000; // 0x2464
	13'h1233: q2 = 16'h3d18; // 0x2466
	13'h1234: q2 = 16'h5c4f; // 0x2468
	13'h1235: q2 = 16'h6032; // 0x246a
	13'h1236: q2 = 16'h7807; // 0x246c
	13'h1237: q2 = 16'h4a44; // 0x246e
	13'h1238: q2 = 16'h6d2c; // 0x2470
	13'h1239: q2 = 16'h3ebc; // 0x2472
	13'h123a: q2 = 16'h003e; // 0x2474
	13'h123b: q2 = 16'h3004; // 0x2476
	13'h123c: q2 = 16'he340; // 0x2478
	13'h123d: q2 = 16'h48c0; // 0x247a
	13'h123e: q2 = 16'hd0bc; // 0x247c
	13'h123f: q2 = 16'h0001; // 0x247e
	13'h1240: q2 = 16'h805c; // 0x2480
	13'h1241: q2 = 16'h2040; // 0x2482
	13'h1242: q2 = 16'h3f10; // 0x2484
	13'h1243: q2 = 16'h0657; // 0x2486
	13'h1244: q2 = 16'h0030; // 0x2488
	13'h1245: q2 = 16'h3f3c; // 0x248a
	13'h1246: q2 = 16'h0006; // 0x248c
	13'h1247: q2 = 16'h3f03; // 0x248e
	13'h1248: q2 = 16'h4eb9; // 0x2490
	13'h1249: q2 = 16'h0000; // 0x2492
	13'h124a: q2 = 16'h3d18; // 0x2494
	13'h124b: q2 = 16'h5c4f; // 0x2496
	13'h124c: q2 = 16'h5543; // 0x2498
	13'h124d: q2 = 16'h5344; // 0x249a
	13'h124e: q2 = 16'h60d0; // 0x249c
	13'h124f: q2 = 16'h5247; // 0x249e
	13'h1250: q2 = 16'h6000; // 0x24a0
	13'h1251: q2 = 16'hfe58; // 0x24a2
	13'h1252: q2 = 16'h526e; // 0x24a4
	13'h1253: q2 = 16'hfffe; // 0x24a6
	13'h1254: q2 = 16'h0c6e; // 0x24a8
	13'h1255: q2 = 16'h000a; // 0x24aa
	13'h1256: q2 = 16'hfffe; // 0x24ac
	13'h1257: q2 = 16'h6612; // 0x24ae
	13'h1258: q2 = 16'h4a79; // 0x24b0
	13'h1259: q2 = 16'h0001; // 0x24b2
	13'h125a: q2 = 16'h758e; // 0x24b4
	13'h125b: q2 = 16'h670a; // 0x24b6
	13'h125c: q2 = 16'h7001; // 0x24b8
	13'h125d: q2 = 16'h9055; // 0x24ba
	13'h125e: q2 = 16'h3a80; // 0x24bc
	13'h125f: q2 = 16'h426e; // 0x24be
	13'h1260: q2 = 16'hfffe; // 0x24c0
	13'h1261: q2 = 16'h4a79; // 0x24c2
	13'h1262: q2 = 16'h0001; // 0x24c4
	13'h1263: q2 = 16'h8a7e; // 0x24c6
	13'h1264: q2 = 16'h670c; // 0x24c8
	13'h1265: q2 = 16'h4a79; // 0x24ca
	13'h1266: q2 = 16'h0001; // 0x24cc
	13'h1267: q2 = 16'h8a80; // 0x24ce
	13'h1268: q2 = 16'h6704; // 0x24d0
	13'h1269: q2 = 16'h4255; // 0x24d2
	13'h126a: q2 = 16'h6004; // 0x24d4
	13'h126b: q2 = 16'h6000; // 0x24d6
	13'h126c: q2 = 16'hfe1a; // 0x24d8
	13'h126d: q2 = 16'h4a9f; // 0x24da
	13'h126e: q2 = 16'h4cdf; // 0x24dc
	13'h126f: q2 = 16'h30f8; // 0x24de
	13'h1270: q2 = 16'h4e5e; // 0x24e0
	13'h1271: q2 = 16'h4e75; // 0x24e2
	13'h1272: q2 = 16'h4e56; // 0x24e4
	13'h1273: q2 = 16'hffdc; // 0x24e6
	13'h1274: q2 = 16'h48e7; // 0x24e8
	13'h1275: q2 = 16'h3f00; // 0x24ea
	13'h1276: q2 = 16'h4246; // 0x24ec
	13'h1277: q2 = 16'h7a01; // 0x24ee
	13'h1278: q2 = 16'h3d7c; // 0x24f0
	13'h1279: q2 = 16'h0001; // 0x24f2
	13'h127a: q2 = 16'hfffe; // 0x24f4
	13'h127b: q2 = 16'h4eb9; // 0x24f6
	13'h127c: q2 = 16'h0000; // 0x24f8
	13'h127d: q2 = 16'h0226; // 0x24fa
	13'h127e: q2 = 16'h4247; // 0x24fc
	13'h127f: q2 = 16'hbe7c; // 0x24fe
	13'h1280: q2 = 16'h0006; // 0x2500
	13'h1281: q2 = 16'h6e60; // 0x2502
	13'h1282: q2 = 16'hbe46; // 0x2504
	13'h1283: q2 = 16'h6604; // 0x2506
	13'h1284: q2 = 16'h762d; // 0x2508
	13'h1285: q2 = 16'h6002; // 0x250a
	13'h1286: q2 = 16'h7636; // 0x250c
	13'h1287: q2 = 16'hbe7c; // 0x250e
	13'h1288: q2 = 16'h0004; // 0x2510
	13'h1289: q2 = 16'h6e04; // 0x2512
	13'h128a: q2 = 16'h7806; // 0x2514
	13'h128b: q2 = 16'h6002; // 0x2516
	13'h128c: q2 = 16'h7864; // 0x2518
	13'h128d: q2 = 16'h3eb9; // 0x251a
	13'h128e: q2 = 16'h0000; // 0x251c
	13'h128f: q2 = 16'hf9be; // 0x251e
	13'h1290: q2 = 16'h3007; // 0x2520
	13'h1291: q2 = 16'hd157; // 0x2522
	13'h1292: q2 = 16'h200e; // 0x2524
	13'h1293: q2 = 16'hd0bc; // 0x2526
	13'h1294: q2 = 16'hffff; // 0x2528
	13'h1295: q2 = 16'hffdc; // 0x252a
	13'h1296: q2 = 16'h2f00; // 0x252c
	13'h1297: q2 = 16'h4eb9; // 0x252e
	13'h1298: q2 = 16'h0000; // 0x2530
	13'h1299: q2 = 16'h78f6; // 0x2532
	13'h129a: q2 = 16'h4a9f; // 0x2534
	13'h129b: q2 = 16'h3e83; // 0x2536
	13'h129c: q2 = 16'h4267; // 0x2538
	13'h129d: q2 = 16'h3f04; // 0x253a
	13'h129e: q2 = 16'h3007; // 0x253c
	13'h129f: q2 = 16'he340; // 0x253e
	13'h12a0: q2 = 16'h48c0; // 0x2540
	13'h12a1: q2 = 16'hd0bc; // 0x2542
	13'h12a2: q2 = 16'h0000; // 0x2544
	13'h12a3: q2 = 16'hf9c0; // 0x2546
	13'h12a4: q2 = 16'h2040; // 0x2548
	13'h12a5: q2 = 16'h3f10; // 0x254a
	13'h12a6: q2 = 16'h200e; // 0x254c
	13'h12a7: q2 = 16'hd0bc; // 0x254e
	13'h12a8: q2 = 16'hffff; // 0x2550
	13'h12a9: q2 = 16'hffdc; // 0x2552
	13'h12aa: q2 = 16'h2f00; // 0x2554
	13'h12ab: q2 = 16'h4eb9; // 0x2556
	13'h12ac: q2 = 16'h0000; // 0x2558
	13'h12ad: q2 = 16'h026c; // 0x255a
	13'h12ae: q2 = 16'hdefc; // 0x255c
	13'h12af: q2 = 16'h000a; // 0x255e
	13'h12b0: q2 = 16'h5247; // 0x2560
	13'h12b1: q2 = 16'h609a; // 0x2562
	13'h12b2: q2 = 16'h3ebc; // 0x2564
	13'h12b3: q2 = 16'h0004; // 0x2566
	13'h12b4: q2 = 16'h3f06; // 0x2568
	13'h12b5: q2 = 16'h4eb9; // 0x256a
	13'h12b6: q2 = 16'h0000; // 0x256c
	13'h12b7: q2 = 16'ha602; // 0x256e
	13'h12b8: q2 = 16'h4a5f; // 0x2570
	13'h12b9: q2 = 16'h3c00; // 0x2572
	13'h12ba: q2 = 16'h4a45; // 0x2574
	13'h12bb: q2 = 16'h6658; // 0x2576
	13'h12bc: q2 = 16'h4a79; // 0x2578
	13'h12bd: q2 = 16'h0001; // 0x257a
	13'h12be: q2 = 16'h7fca; // 0x257c
	13'h12bf: q2 = 16'h6750; // 0x257e
	13'h12c0: q2 = 16'h3006; // 0x2580
	13'h12c1: q2 = 16'h602a; // 0x2582
	13'h12c2: q2 = 16'h4eb9; // 0x2584
	13'h12c3: q2 = 16'h0000; // 0x2586
	13'h12c4: q2 = 16'h9b50; // 0x2588
	13'h12c5: q2 = 16'h6036; // 0x258a
	13'h12c6: q2 = 16'h4eb9; // 0x258c
	13'h12c7: q2 = 16'h0000; // 0x258e
	13'h12c8: q2 = 16'ha258; // 0x2590
	13'h12c9: q2 = 16'h602e; // 0x2592
	13'h12ca: q2 = 16'h4eb9; // 0x2594
	13'h12cb: q2 = 16'h0000; // 0x2596
	13'h12cc: q2 = 16'h99fe; // 0x2598
	13'h12cd: q2 = 16'h6026; // 0x259a
	13'h12ce: q2 = 16'h4eb9; // 0x259c
	13'h12cf: q2 = 16'h0000; // 0x259e
	13'h12d0: q2 = 16'h9ae4; // 0x25a0
	13'h12d1: q2 = 16'h601e; // 0x25a2
	13'h12d2: q2 = 16'h4eb9; // 0x25a4
	13'h12d3: q2 = 16'h0000; // 0x25a6
	13'h12d4: q2 = 16'ha136; // 0x25a8
	13'h12d5: q2 = 16'h6016; // 0x25aa
	13'h12d6: q2 = 16'h6014; // 0x25ac
	13'h12d7: q2 = 16'hb07c; // 0x25ae
	13'h12d8: q2 = 16'h0004; // 0x25b0
	13'h12d9: q2 = 16'h620e; // 0x25b2
	13'h12da: q2 = 16'he540; // 0x25b4
	13'h12db: q2 = 16'h3040; // 0x25b6
	13'h12dc: q2 = 16'hd1fc; // 0x25b8
	13'h12dd: q2 = 16'h0000; // 0x25ba
	13'h12de: q2 = 16'hfabe; // 0x25bc
	13'h12df: q2 = 16'h2050; // 0x25be
	13'h12e0: q2 = 16'h4ed0; // 0x25c0
	13'h12e1: q2 = 16'h4eb9; // 0x25c2
	13'h12e2: q2 = 16'h0000; // 0x25c4
	13'h12e3: q2 = 16'h0226; // 0x25c6
	13'h12e4: q2 = 16'h7a01; // 0x25c8
	13'h12e5: q2 = 16'h3d7c; // 0x25ca
	13'h12e6: q2 = 16'h0001; // 0x25cc
	13'h12e7: q2 = 16'hfffe; // 0x25ce
	13'h12e8: q2 = 16'h4a79; // 0x25d0
	13'h12e9: q2 = 16'h0001; // 0x25d2
	13'h12ea: q2 = 16'h7fca; // 0x25d4
	13'h12eb: q2 = 16'h6602; // 0x25d6
	13'h12ec: q2 = 16'h4245; // 0x25d8
	13'h12ed: q2 = 16'h4a79; // 0x25da
	13'h12ee: q2 = 16'h0001; // 0x25dc
	13'h12ef: q2 = 16'h8a7e; // 0x25de
	13'h12f0: q2 = 16'h6604; // 0x25e0
	13'h12f1: q2 = 16'h426e; // 0x25e2
	13'h12f2: q2 = 16'hfffe; // 0x25e4
	13'h12f3: q2 = 16'h4a6e; // 0x25e6
	13'h12f4: q2 = 16'hfffe; // 0x25e8
	13'h12f5: q2 = 16'h6608; // 0x25ea
	13'h12f6: q2 = 16'h4a79; // 0x25ec
	13'h12f7: q2 = 16'h0001; // 0x25ee
	13'h12f8: q2 = 16'h8a7e; // 0x25f0
	13'h12f9: q2 = 16'h6604; // 0x25f2
	13'h12fa: q2 = 16'h6000; // 0x25f4
	13'h12fb: q2 = 16'hff06; // 0x25f6
	13'h12fc: q2 = 16'h4a9f; // 0x25f8
	13'h12fd: q2 = 16'h4cdf; // 0x25fa
	13'h12fe: q2 = 16'h00f8; // 0x25fc
	13'h12ff: q2 = 16'h4e5e; // 0x25fe
	13'h1300: q2 = 16'h4e75; // 0x2600
	13'h1301: q2 = 16'h4e56; // 0x2602
	13'h1302: q2 = 16'h0000; // 0x2604
	13'h1303: q2 = 16'h48e7; // 0x2606
	13'h1304: q2 = 16'h0700; // 0x2608
	13'h1305: q2 = 16'h3e2e; // 0x260a
	13'h1306: q2 = 16'h0008; // 0x260c
	13'h1307: q2 = 16'h3c2e; // 0x260e
	13'h1308: q2 = 16'h000a; // 0x2610
	13'h1309: q2 = 16'h4a79; // 0x2612
	13'h130a: q2 = 16'h0001; // 0x2614
	13'h130b: q2 = 16'h7fca; // 0x2616
	13'h130c: q2 = 16'h6600; // 0x2618
	13'h130d: q2 = 16'h010a; // 0x261a
	13'h130e: q2 = 16'h4ab9; // 0x261c
	13'h130f: q2 = 16'h0001; // 0x261e
	13'h1310: q2 = 16'h7fc2; // 0x2620
	13'h1311: q2 = 16'h6600; // 0x2622
	13'h1312: q2 = 16'h0076; // 0x2624
	13'h1313: q2 = 16'h4a79; // 0x2626
	13'h1314: q2 = 16'h0001; // 0x2628
	13'h1315: q2 = 16'h8a80; // 0x262a
	13'h1316: q2 = 16'h666c; // 0x262c
	13'h1317: q2 = 16'h2079; // 0x262e
	13'h1318: q2 = 16'h0001; // 0x2630
	13'h1319: q2 = 16'h7eb2; // 0x2632
	13'h131a: q2 = 16'h3028; // 0x2634
	13'h131b: q2 = 16'h0004; // 0x2636
	13'h131c: q2 = 16'h2279; // 0x2638
	13'h131d: q2 = 16'h0001; // 0x263a
	13'h131e: q2 = 16'h7eb2; // 0x263c
	13'h131f: q2 = 16'h9069; // 0x263e
	13'h1320: q2 = 16'h0006; // 0x2640
	13'h1321: q2 = 16'he440; // 0x2642
	13'h1322: q2 = 16'hb079; // 0x2644
	13'h1323: q2 = 16'h0001; // 0x2646
	13'h1324: q2 = 16'h8624; // 0x2648
	13'h1325: q2 = 16'h6f14; // 0x264a
	13'h1326: q2 = 16'h5247; // 0x264c
	13'h1327: q2 = 16'hbe46; // 0x264e
	13'h1328: q2 = 16'h6f02; // 0x2650
	13'h1329: q2 = 16'h4247; // 0x2652
	13'h132a: q2 = 16'h23fc; // 0x2654
	13'h132b: q2 = 16'h0000; // 0x2656
	13'h132c: q2 = 16'h0012; // 0x2658
	13'h132d: q2 = 16'h0001; // 0x265a
	13'h132e: q2 = 16'h7fc2; // 0x265c
	13'h132f: q2 = 16'h6030; // 0x265e
	13'h1330: q2 = 16'h2079; // 0x2660
	13'h1331: q2 = 16'h0001; // 0x2662
	13'h1332: q2 = 16'h7eb2; // 0x2664
	13'h1333: q2 = 16'h3028; // 0x2666
	13'h1334: q2 = 16'h0006; // 0x2668
	13'h1335: q2 = 16'h2279; // 0x266a
	13'h1336: q2 = 16'h0001; // 0x266c
	13'h1337: q2 = 16'h7eb2; // 0x266e
	13'h1338: q2 = 16'h9069; // 0x2670
	13'h1339: q2 = 16'h0004; // 0x2672
	13'h133a: q2 = 16'he440; // 0x2674
	13'h133b: q2 = 16'hb079; // 0x2676
	13'h133c: q2 = 16'h0001; // 0x2678
	13'h133d: q2 = 16'h8624; // 0x267a
	13'h133e: q2 = 16'h6c12; // 0x267c
	13'h133f: q2 = 16'h5347; // 0x267e
	13'h1340: q2 = 16'h4a47; // 0x2680
	13'h1341: q2 = 16'h6c02; // 0x2682
	13'h1342: q2 = 16'h3e06; // 0x2684
	13'h1343: q2 = 16'h23fc; // 0x2686
	13'h1344: q2 = 16'h0000; // 0x2688
	13'h1345: q2 = 16'h0012; // 0x268a
	13'h1346: q2 = 16'h0001; // 0x268c
	13'h1347: q2 = 16'h7fc2; // 0x268e
	13'h1348: q2 = 16'h4279; // 0x2690
	13'h1349: q2 = 16'h0001; // 0x2692
	13'h134a: q2 = 16'h85fc; // 0x2694
	13'h134b: q2 = 16'h6000; // 0x2696
	13'h134c: q2 = 16'h008c; // 0x2698
	13'h134d: q2 = 16'h4a79; // 0x269a
	13'h134e: q2 = 16'h0001; // 0x269c
	13'h134f: q2 = 16'h8a80; // 0x269e
	13'h1350: q2 = 16'h6714; // 0x26a0
	13'h1351: q2 = 16'h4a79; // 0x26a2
	13'h1352: q2 = 16'h0001; // 0x26a4
	13'h1353: q2 = 16'h85fc; // 0x26a6
	13'h1354: q2 = 16'h660c; // 0x26a8
	13'h1355: q2 = 16'h33fc; // 0x26aa
	13'h1356: q2 = 16'h0001; // 0x26ac
	13'h1357: q2 = 16'h0001; // 0x26ae
	13'h1358: q2 = 16'h85fc; // 0x26b0
	13'h1359: q2 = 16'h6000; // 0x26b2
	13'h135a: q2 = 16'h0070; // 0x26b4
	13'h135b: q2 = 16'h4a79; // 0x26b6
	13'h135c: q2 = 16'h0001; // 0x26b8
	13'h135d: q2 = 16'h8a80; // 0x26ba
	13'h135e: q2 = 16'h6716; // 0x26bc
	13'h135f: q2 = 16'h0c79; // 0x26be
	13'h1360: q2 = 16'h0001; // 0x26c0
	13'h1361: q2 = 16'h0001; // 0x26c2
	13'h1362: q2 = 16'h85fc; // 0x26c4
	13'h1363: q2 = 16'h660c; // 0x26c6
	13'h1364: q2 = 16'h23fc; // 0x26c8
	13'h1365: q2 = 16'h0000; // 0x26ca
	13'h1366: q2 = 16'h0012; // 0x26cc
	13'h1367: q2 = 16'h0001; // 0x26ce
	13'h1368: q2 = 16'h7fc2; // 0x26d0
	13'h1369: q2 = 16'h6050; // 0x26d2
	13'h136a: q2 = 16'h4a79; // 0x26d4
	13'h136b: q2 = 16'h0001; // 0x26d6
	13'h136c: q2 = 16'h8a80; // 0x26d8
	13'h136d: q2 = 16'h6726; // 0x26da
	13'h136e: q2 = 16'h0c79; // 0x26dc
	13'h136f: q2 = 16'h0002; // 0x26de
	13'h1370: q2 = 16'h0001; // 0x26e0
	13'h1371: q2 = 16'h85fc; // 0x26e2
	13'h1372: q2 = 16'h661c; // 0x26e4
	13'h1373: q2 = 16'h33fc; // 0x26e6
	13'h1374: q2 = 16'h0001; // 0x26e8
	13'h1375: q2 = 16'h0001; // 0x26ea
	13'h1376: q2 = 16'h85fc; // 0x26ec
	13'h1377: q2 = 16'h5247; // 0x26ee
	13'h1378: q2 = 16'hbe46; // 0x26f0
	13'h1379: q2 = 16'h6f02; // 0x26f2
	13'h137a: q2 = 16'h4247; // 0x26f4
	13'h137b: q2 = 16'h23fc; // 0x26f6
	13'h137c: q2 = 16'h0000; // 0x26f8
	13'h137d: q2 = 16'h0012; // 0x26fa
	13'h137e: q2 = 16'h0001; // 0x26fc
	13'h137f: q2 = 16'h7fc2; // 0x26fe
	13'h1380: q2 = 16'h6022; // 0x2700
	13'h1381: q2 = 16'h4ab9; // 0x2702
	13'h1382: q2 = 16'h0001; // 0x2704
	13'h1383: q2 = 16'h7fc2; // 0x2706
	13'h1384: q2 = 16'h671a; // 0x2708
	13'h1385: q2 = 16'h4a79; // 0x270a
	13'h1386: q2 = 16'h0001; // 0x270c
	13'h1387: q2 = 16'h8a80; // 0x270e
	13'h1388: q2 = 16'h6612; // 0x2710
	13'h1389: q2 = 16'h0c79; // 0x2712
	13'h138a: q2 = 16'h0001; // 0x2714
	13'h138b: q2 = 16'h0001; // 0x2716
	13'h138c: q2 = 16'h85fc; // 0x2718
	13'h138d: q2 = 16'h6608; // 0x271a
	13'h138e: q2 = 16'h33fc; // 0x271c
	13'h138f: q2 = 16'h0002; // 0x271e
	13'h1390: q2 = 16'h0001; // 0x2720
	13'h1391: q2 = 16'h85fc; // 0x2722
	13'h1392: q2 = 16'h3007; // 0x2724
	13'h1393: q2 = 16'h4a9f; // 0x2726
	13'h1394: q2 = 16'h4cdf; // 0x2728
	13'h1395: q2 = 16'h00c0; // 0x272a
	13'h1396: q2 = 16'h4e5e; // 0x272c
	13'h1397: q2 = 16'h4e75; // 0x272e
	13'h1398: q2 = 16'h4e56; // 0x2730
	13'h1399: q2 = 16'h0000; // 0x2732
	13'h139a: q2 = 16'h48e7; // 0x2734
	13'h139b: q2 = 16'h3f00; // 0x2736
	13'h139c: q2 = 16'h3e2e; // 0x2738
	13'h139d: q2 = 16'h000a; // 0x273a
	13'h139e: q2 = 16'h3a2e; // 0x273c
	13'h139f: q2 = 16'h0008; // 0x273e
	13'h13a0: q2 = 16'h4244; // 0x2740
	13'h13a1: q2 = 16'hba7c; // 0x2742
	13'h13a2: q2 = 16'h0023; // 0x2744
	13'h13a3: q2 = 16'h6f06; // 0x2746
	13'h13a4: q2 = 16'h7801; // 0x2748
	13'h13a5: q2 = 16'h9a7c; // 0x274a
	13'h13a6: q2 = 16'h0024; // 0x274c
	13'h13a7: q2 = 16'h3005; // 0x274e
	13'h13a8: q2 = 16'h48c0; // 0x2750
	13'h13a9: q2 = 16'hd0bc; // 0x2752
	13'h13aa: q2 = 16'h0000; // 0x2754
	13'h13ab: q2 = 16'hfad2; // 0x2756
	13'h13ac: q2 = 16'h2040; // 0x2758
	13'h13ad: q2 = 16'h1c10; // 0x275a
	13'h13ae: q2 = 16'h4886; // 0x275c
	13'h13af: q2 = 16'hcc7c; // 0x275e
	13'h13b0: q2 = 16'h00ff; // 0x2760
	13'h13b1: q2 = 16'hba7c; // 0x2762
	13'h13b2: q2 = 16'h0012; // 0x2764
	13'h13b3: q2 = 16'h6604; // 0x2766
	13'h13b4: q2 = 16'h3c3c; // 0x2768
	13'h13b5: q2 = 16'h0100; // 0x276a
	13'h13b6: q2 = 16'h3006; // 0x276c
	13'h13b7: q2 = 16'hc1c7; // 0x276e
	13'h13b8: q2 = 16'h2600; // 0x2770
	13'h13b9: q2 = 16'h2003; // 0x2772
	13'h13ba: q2 = 16'he080; // 0x2774
	13'h13bb: q2 = 16'h2600; // 0x2776
	13'h13bc: q2 = 16'h2003; // 0x2778
	13'h13bd: q2 = 16'h3c00; // 0x277a
	13'h13be: q2 = 16'h4a44; // 0x277c
	13'h13bf: q2 = 16'h6706; // 0x277e
	13'h13c0: q2 = 16'h3006; // 0x2780
	13'h13c1: q2 = 16'h4440; // 0x2782
	13'h13c2: q2 = 16'h3c00; // 0x2784
	13'h13c3: q2 = 16'h3006; // 0x2786
	13'h13c4: q2 = 16'h4a9f; // 0x2788
	13'h13c5: q2 = 16'h4cdf; // 0x278a
	13'h13c6: q2 = 16'h00f8; // 0x278c
	13'h13c7: q2 = 16'h4e5e; // 0x278e
	13'h13c8: q2 = 16'h4e75; // 0x2790
	13'h13c9: q2 = 16'h4e56; // 0x2792
	13'h13ca: q2 = 16'hfff4; // 0x2794
	13'h13cb: q2 = 16'h48e7; // 0x2796
	13'h13cc: q2 = 16'h3f0c; // 0x2798
	13'h13cd: q2 = 16'h33fc; // 0x279a
	13'h13ce: q2 = 16'h0001; // 0x279c
	13'h13cf: q2 = 16'h0001; // 0x279e
	13'h13d0: q2 = 16'h7f2a; // 0x27a0
	13'h13d1: q2 = 16'h4eb9; // 0x27a2
	13'h13d2: q2 = 16'h0000; // 0x27a4
	13'h13d3: q2 = 16'h4ee2; // 0x27a6
	13'h13d4: q2 = 16'h3c00; // 0x27a8
	13'h13d5: q2 = 16'h4eb9; // 0x27aa
	13'h13d6: q2 = 16'h0000; // 0x27ac
	13'h13d7: q2 = 16'h4f30; // 0x27ae
	13'h13d8: q2 = 16'h3a00; // 0x27b0
	13'h13d9: q2 = 16'h426e; // 0x27b2
	13'h13da: q2 = 16'hfff4; // 0x27b4
	13'h13db: q2 = 16'h287c; // 0x27b6
	13'h13dc: q2 = 16'h0001; // 0x27b8
	13'h13dd: q2 = 16'h893e; // 0x27ba
	13'h13de: q2 = 16'h4247; // 0x27bc
	13'h13df: q2 = 16'hbe79; // 0x27be
	13'h13e0: q2 = 16'h0001; // 0x27c0
	13'h13e1: q2 = 16'h7fa8; // 0x27c2
	13'h13e2: q2 = 16'h6c1a; // 0x27c4
	13'h13e3: q2 = 16'h0c6c; // 0x27c6
	13'h13e4: q2 = 16'h0005; // 0x27c8
	13'h13e5: q2 = 16'h0004; // 0x27ca
	13'h13e6: q2 = 16'h6708; // 0x27cc
	13'h13e7: q2 = 16'h302c; // 0x27ce
	13'h13e8: q2 = 16'h0006; // 0x27d0
	13'h13e9: q2 = 16'hd16e; // 0x27d2
	13'h13ea: q2 = 16'hfff4; // 0x27d4
	13'h13eb: q2 = 16'hd9fc; // 0x27d6
	13'h13ec: q2 = 16'h0000; // 0x27d8
	13'h13ed: q2 = 16'h0010; // 0x27da
	13'h13ee: q2 = 16'h5247; // 0x27dc
	13'h13ef: q2 = 16'h60de; // 0x27de
	13'h13f0: q2 = 16'h426e; // 0x27e0
	13'h13f1: q2 = 16'hfff8; // 0x27e2
	13'h13f2: q2 = 16'h23fc; // 0x27e4
	13'h13f3: q2 = 16'h0000; // 0x27e6
	13'h13f4: q2 = 16'h0002; // 0x27e8
	13'h13f5: q2 = 16'h0001; // 0x27ea
	13'h13f6: q2 = 16'h7fc2; // 0x27ec
	13'h13f7: q2 = 16'h287c; // 0x27ee
	13'h13f8: q2 = 16'h0001; // 0x27f0
	13'h13f9: q2 = 16'h893e; // 0x27f2
	13'h13fa: q2 = 16'h4247; // 0x27f4
	13'h13fb: q2 = 16'hbe79; // 0x27f6
	13'h13fc: q2 = 16'h0001; // 0x27f8
	13'h13fd: q2 = 16'h7fa8; // 0x27fa
	13'h13fe: q2 = 16'h6c00; // 0x27fc
	13'h13ff: q2 = 16'h0132; // 0x27fe
	13'h1400: q2 = 16'h0c6e; // 0x2800
	13'h1401: q2 = 16'h001a; // 0x2802
	13'h1402: q2 = 16'hfff8; // 0x2804
	13'h1403: q2 = 16'h6f08; // 0x2806
	13'h1404: q2 = 16'h4a6e; // 0x2808
	13'h1405: q2 = 16'hfff4; // 0x280a
	13'h1406: q2 = 16'h6700; // 0x280c
	13'h1407: q2 = 16'h0122; // 0x280e
	13'h1408: q2 = 16'h0c6c; // 0x2810
	13'h1409: q2 = 16'h0005; // 0x2812
	13'h140a: q2 = 16'h0004; // 0x2814
	13'h140b: q2 = 16'h6708; // 0x2816
	13'h140c: q2 = 16'h4a6c; // 0x2818
	13'h140d: q2 = 16'h0006; // 0x281a
	13'h140e: q2 = 16'h6600; // 0x281c
	13'h140f: q2 = 16'h007e; // 0x281e
	13'h1410: q2 = 16'h3ebc; // 0x2820
	13'h1411: q2 = 16'h7880; // 0x2822
	13'h1412: q2 = 16'h3f3c; // 0x2824
	13'h1413: q2 = 16'h0080; // 0x2826
	13'h1414: q2 = 16'h4eb9; // 0x2828
	13'h1415: q2 = 16'h0000; // 0x282a
	13'h1416: q2 = 16'h8e6c; // 0x282c
	13'h1417: q2 = 16'h4a5f; // 0x282e
	13'h1418: q2 = 16'h3800; // 0x2830
	13'h1419: q2 = 16'h3ebc; // 0x2832
	13'h141a: q2 = 16'h7800; // 0x2834
	13'h141b: q2 = 16'h3f3c; // 0x2836
	13'h141c: q2 = 16'h1280; // 0x2838
	13'h141d: q2 = 16'h4eb9; // 0x283a
	13'h141e: q2 = 16'h0000; // 0x283c
	13'h141f: q2 = 16'h8e6c; // 0x283e
	13'h1420: q2 = 16'h4a5f; // 0x2840
	13'h1421: q2 = 16'h3600; // 0x2842
	13'h1422: q2 = 16'h3ebc; // 0x2844
	13'h1423: q2 = 16'h0003; // 0x2846
	13'h1424: q2 = 16'h4267; // 0x2848
	13'h1425: q2 = 16'h4eb9; // 0x284a
	13'h1426: q2 = 16'h0000; // 0x284c
	13'h1427: q2 = 16'h8e6c; // 0x284e
	13'h1428: q2 = 16'h4a5f; // 0x2850
	13'h1429: q2 = 16'h3d40; // 0x2852
	13'h142a: q2 = 16'hfff6; // 0x2854
	13'h142b: q2 = 16'h4a6e; // 0x2856
	13'h142c: q2 = 16'hfff6; // 0x2858
	13'h142d: q2 = 16'h6606; // 0x285a
	13'h142e: q2 = 16'h383c; // 0x285c
	13'h142f: q2 = 16'h0080; // 0x285e
	13'h1430: q2 = 16'h6028; // 0x2860
	13'h1431: q2 = 16'h0c6e; // 0x2862
	13'h1432: q2 = 16'h0001; // 0x2864
	13'h1433: q2 = 16'hfff6; // 0x2866
	13'h1434: q2 = 16'h6606; // 0x2868
	13'h1435: q2 = 16'h383c; // 0x286a
	13'h1436: q2 = 16'h7880; // 0x286c
	13'h1437: q2 = 16'h601a; // 0x286e
	13'h1438: q2 = 16'h0c6e; // 0x2870
	13'h1439: q2 = 16'h0002; // 0x2872
	13'h143a: q2 = 16'hfff6; // 0x2874
	13'h143b: q2 = 16'h6606; // 0x2876
	13'h143c: q2 = 16'h363c; // 0x2878
	13'h143d: q2 = 16'h1280; // 0x287a
	13'h143e: q2 = 16'h600c; // 0x287c
	13'h143f: q2 = 16'h0c6e; // 0x287e
	13'h1440: q2 = 16'h0003; // 0x2880
	13'h1441: q2 = 16'hfff6; // 0x2882
	13'h1442: q2 = 16'h6604; // 0x2884
	13'h1443: q2 = 16'h363c; // 0x2886
	13'h1444: q2 = 16'h7800; // 0x2888
	13'h1445: q2 = 16'h3eb9; // 0x288a
	13'h1446: q2 = 16'h0001; // 0x288c
	13'h1447: q2 = 16'h8070; // 0x288e
	13'h1448: q2 = 16'h4eb9; // 0x2890
	13'h1449: q2 = 16'h0000; // 0x2892
	13'h144a: q2 = 16'h3e52; // 0x2894
	13'h144b: q2 = 16'h3d40; // 0x2896
	13'h144c: q2 = 16'hfffa; // 0x2898
	13'h144d: q2 = 16'h6026; // 0x289a
	13'h144e: q2 = 16'h382c; // 0x289c
	13'h144f: q2 = 16'h0008; // 0x289e
	13'h1450: q2 = 16'h362c; // 0x28a0
	13'h1451: q2 = 16'h000a; // 0x28a2
	13'h1452: q2 = 16'h3d6c; // 0x28a4
	13'h1453: q2 = 16'h0004; // 0x28a6
	13'h1454: q2 = 16'hfffa; // 0x28a8
	13'h1455: q2 = 16'h536c; // 0x28aa
	13'h1456: q2 = 16'h0006; // 0x28ac
	13'h1457: q2 = 16'h2e8c; // 0x28ae
	13'h1458: q2 = 16'h4eb9; // 0x28b0
	13'h1459: q2 = 16'h0000; // 0x28b2
	13'h145a: q2 = 16'h161a; // 0x28b4
	13'h145b: q2 = 16'h2e8c; // 0x28b6
	13'h145c: q2 = 16'h4eb9; // 0x28b8
	13'h145d: q2 = 16'h0000; // 0x28ba
	13'h145e: q2 = 16'h0f60; // 0x28bc
	13'h145f: q2 = 16'h536e; // 0x28be
	13'h1460: q2 = 16'hfff4; // 0x28c0
	13'h1461: q2 = 16'h3e83; // 0x28c2
	13'h1462: q2 = 16'h3f04; // 0x28c4
	13'h1463: q2 = 16'h3f2e; // 0x28c6
	13'h1464: q2 = 16'hfffa; // 0x28c8
	13'h1465: q2 = 16'h4eb9; // 0x28ca
	13'h1466: q2 = 16'h0000; // 0x28cc
	13'h1467: q2 = 16'h38d8; // 0x28ce
	13'h1468: q2 = 16'h4a9f; // 0x28d0
	13'h1469: q2 = 16'h2a40; // 0x28d2
	13'h146a: q2 = 16'h200d; // 0x28d4
	13'h146b: q2 = 16'h674c; // 0x28d6
	13'h146c: q2 = 16'h3006; // 0x28d8
	13'h146d: q2 = 16'h9044; // 0x28da
	13'h146e: q2 = 16'h3d40; // 0x28dc
	13'h146f: q2 = 16'hfffe; // 0x28de
	13'h1470: q2 = 16'h3005; // 0x28e0
	13'h1471: q2 = 16'h9043; // 0x28e2
	13'h1472: q2 = 16'h3d40; // 0x28e4
	13'h1473: q2 = 16'hfffc; // 0x28e6
	13'h1474: q2 = 16'h200e; // 0x28e8
	13'h1475: q2 = 16'hd0bc; // 0x28ea
	13'h1476: q2 = 16'hffff; // 0x28ec
	13'h1477: q2 = 16'hfffc; // 0x28ee
	13'h1478: q2 = 16'h2e80; // 0x28f0
	13'h1479: q2 = 16'h200e; // 0x28f2
	13'h147a: q2 = 16'hd0bc; // 0x28f4
	13'h147b: q2 = 16'hffff; // 0x28f6
	13'h147c: q2 = 16'hfffe; // 0x28f8
	13'h147d: q2 = 16'h2f00; // 0x28fa
	13'h147e: q2 = 16'h3f3c; // 0x28fc
	13'h147f: q2 = 16'h0400; // 0x28fe
	13'h1480: q2 = 16'h4eb9; // 0x2900
	13'h1481: q2 = 16'h0000; // 0x2902
	13'h1482: q2 = 16'h09bc; // 0x2904
	13'h1483: q2 = 16'h5c4f; // 0x2906
	13'h1484: q2 = 16'h3e85; // 0x2908
	13'h1485: q2 = 16'h3f06; // 0x290a
	13'h1486: q2 = 16'h3f2e; // 0x290c
	13'h1487: q2 = 16'hfffc; // 0x290e
	13'h1488: q2 = 16'h3f2e; // 0x2910
	13'h1489: q2 = 16'hfffe; // 0x2912
	13'h148a: q2 = 16'h2f0d; // 0x2914
	13'h148b: q2 = 16'h4eb9; // 0x2916
	13'h148c: q2 = 16'h0000; // 0x2918
	13'h148d: q2 = 16'h3988; // 0x291a
	13'h148e: q2 = 16'hdefc; // 0x291c
	13'h148f: q2 = 16'h000a; // 0x291e
	13'h1490: q2 = 16'h526e; // 0x2920
	13'h1491: q2 = 16'hfff8; // 0x2922
	13'h1492: q2 = 16'hd9fc; // 0x2924
	13'h1493: q2 = 16'h0000; // 0x2926
	13'h1494: q2 = 16'h0010; // 0x2928
	13'h1495: q2 = 16'h5247; // 0x292a
	13'h1496: q2 = 16'h6000; // 0x292c
	13'h1497: q2 = 16'hfec8; // 0x292e
	13'h1498: q2 = 16'h4eb9; // 0x2930
	13'h1499: q2 = 16'h0000; // 0x2932
	13'h149a: q2 = 16'h2fb4; // 0x2934
	13'h149b: q2 = 16'h4eb9; // 0x2936
	13'h149c: q2 = 16'h0000; // 0x2938
	13'h149d: q2 = 16'h18d0; // 0x293a
	13'h149e: q2 = 16'h4eb9; // 0x293c
	13'h149f: q2 = 16'h0000; // 0x293e
	13'h14a0: q2 = 16'h3396; // 0x2940
	13'h14a1: q2 = 16'h4a40; // 0x2942
	13'h14a2: q2 = 16'h660e; // 0x2944
	13'h14a3: q2 = 16'h4ab9; // 0x2946
	13'h14a4: q2 = 16'h0001; // 0x2948
	13'h14a5: q2 = 16'h7fc2; // 0x294a
	13'h14a6: q2 = 16'h6702; // 0x294c
	13'h14a7: q2 = 16'h60f6; // 0x294e
	13'h14a8: q2 = 16'h6000; // 0x2950
	13'h14a9: q2 = 16'hfe92; // 0x2952
	13'h14aa: q2 = 16'h4279; // 0x2954
	13'h14ab: q2 = 16'h0001; // 0x2956
	13'h14ac: q2 = 16'h7f2a; // 0x2958
	13'h14ad: q2 = 16'h4a9f; // 0x295a
	13'h14ae: q2 = 16'h4cdf; // 0x295c
	13'h14af: q2 = 16'h30f8; // 0x295e
	13'h14b0: q2 = 16'h4e5e; // 0x2960
	13'h14b1: q2 = 16'h4e75; // 0x2962
	13'h14b2: q2 = 16'h4e56; // 0x2964
	13'h14b3: q2 = 16'h0000; // 0x2966
	13'h14b4: q2 = 16'h48e7; // 0x2968
	13'h14b5: q2 = 16'h0300; // 0x296a
	13'h14b6: q2 = 16'h23f9; // 0x296c
	13'h14b7: q2 = 16'h0001; // 0x296e
	13'h14b8: q2 = 16'h75ca; // 0x2970
	13'h14b9: q2 = 16'h0001; // 0x2972
	13'h14ba: q2 = 16'h75d6; // 0x2974
	13'h14bb: q2 = 16'h4247; // 0x2976
	13'h14bc: q2 = 16'hbe7c; // 0x2978
	13'h14bd: q2 = 16'h0001; // 0x297a
	13'h14be: q2 = 16'h6e26; // 0x297c
	13'h14bf: q2 = 16'h3007; // 0x297e
	13'h14c0: q2 = 16'he340; // 0x2980
	13'h14c1: q2 = 16'h48c0; // 0x2982
	13'h14c2: q2 = 16'hd0bc; // 0x2984
	13'h14c3: q2 = 16'h0001; // 0x2986
	13'h14c4: q2 = 16'h75da; // 0x2988
	13'h14c5: q2 = 16'h2040; // 0x298a
	13'h14c6: q2 = 16'h4250; // 0x298c
	13'h14c7: q2 = 16'h3007; // 0x298e
	13'h14c8: q2 = 16'he540; // 0x2990
	13'h14c9: q2 = 16'h48c0; // 0x2992
	13'h14ca: q2 = 16'hd0bc; // 0x2994
	13'h14cb: q2 = 16'h0001; // 0x2996
	13'h14cc: q2 = 16'h75de; // 0x2998
	13'h14cd: q2 = 16'h2040; // 0x299a
	13'h14ce: q2 = 16'h7000; // 0x299c
	13'h14cf: q2 = 16'h2080; // 0x299e
	13'h14d0: q2 = 16'h5247; // 0x29a0
	13'h14d1: q2 = 16'h60d4; // 0x29a2
	13'h14d2: q2 = 16'h4a9f; // 0x29a4
	13'h14d3: q2 = 16'h4cdf; // 0x29a6
	13'h14d4: q2 = 16'h0080; // 0x29a8
	13'h14d5: q2 = 16'h4e5e; // 0x29aa
	13'h14d6: q2 = 16'h4e75; // 0x29ac
	13'h14d7: q2 = 16'h4e56; // 0x29ae
	13'h14d8: q2 = 16'h0000; // 0x29b0
	13'h14d9: q2 = 16'h48e7; // 0x29b2
	13'h14da: q2 = 16'h0700; // 0x29b4
	13'h14db: q2 = 16'h3e2e; // 0x29b6
	13'h14dc: q2 = 16'h0008; // 0x29b8
	13'h14dd: q2 = 16'h4a47; // 0x29ba
	13'h14de: q2 = 16'h6610; // 0x29bc
	13'h14df: q2 = 16'h4ab9; // 0x29be
	13'h14e0: q2 = 16'h0001; // 0x29c0
	13'h14e1: q2 = 16'h75e2; // 0x29c2
	13'h14e2: q2 = 16'h6608; // 0x29c4
	13'h14e3: q2 = 16'h52b9; // 0x29c6
	13'h14e4: q2 = 16'h0001; // 0x29c8
	13'h14e5: q2 = 16'h759a; // 0x29ca
	13'h14e6: q2 = 16'h600c; // 0x29cc
	13'h14e7: q2 = 16'hbe7c; // 0x29ce
	13'h14e8: q2 = 16'h0001; // 0x29d0
	13'h14e9: q2 = 16'h6606; // 0x29d2
	13'h14ea: q2 = 16'h52b9; // 0x29d4
	13'h14eb: q2 = 16'h0001; // 0x29d6
	13'h14ec: q2 = 16'h759e; // 0x29d8
	13'h14ed: q2 = 16'h2039; // 0x29da
	13'h14ee: q2 = 16'h0001; // 0x29dc
	13'h14ef: q2 = 16'h75ca; // 0x29de
	13'h14f0: q2 = 16'h90b9; // 0x29e0
	13'h14f1: q2 = 16'h0001; // 0x29e2
	13'h14f2: q2 = 16'h75d6; // 0x29e4
	13'h14f3: q2 = 16'h2f00; // 0x29e6
	13'h14f4: q2 = 16'h3007; // 0x29e8
	13'h14f5: q2 = 16'he540; // 0x29ea
	13'h14f6: q2 = 16'h48c0; // 0x29ec
	13'h14f7: q2 = 16'hd0bc; // 0x29ee
	13'h14f8: q2 = 16'h0001; // 0x29f0
	13'h14f9: q2 = 16'h75de; // 0x29f2
	13'h14fa: q2 = 16'h2040; // 0x29f4
	13'h14fb: q2 = 16'h2010; // 0x29f6
	13'h14fc: q2 = 16'h221f; // 0x29f8
	13'h14fd: q2 = 16'hd081; // 0x29fa
	13'h14fe: q2 = 16'h2c00; // 0x29fc
	13'h14ff: q2 = 16'hddb9; // 0x29fe
	13'h1500: q2 = 16'h0001; // 0x2a00
	13'h1501: q2 = 16'h75c2; // 0x2a02
	13'h1502: q2 = 16'hbcb9; // 0x2a04
	13'h1503: q2 = 16'h0001; // 0x2a06
	13'h1504: q2 = 16'h75c6; // 0x2a08
	13'h1505: q2 = 16'h6f06; // 0x2a0a
	13'h1506: q2 = 16'h23c6; // 0x2a0c
	13'h1507: q2 = 16'h0001; // 0x2a0e
	13'h1508: q2 = 16'h75c6; // 0x2a10
	13'h1509: q2 = 16'h3007; // 0x2a12
	13'h150a: q2 = 16'he340; // 0x2a14
	13'h150b: q2 = 16'h48c0; // 0x2a16
	13'h150c: q2 = 16'hd0bc; // 0x2a18
	13'h150d: q2 = 16'h0001; // 0x2a1a
	13'h150e: q2 = 16'h75da; // 0x2a1c
	13'h150f: q2 = 16'h2040; // 0x2a1e
	13'h1510: q2 = 16'h4a50; // 0x2a20
	13'h1511: q2 = 16'h6f06; // 0x2a22
	13'h1512: q2 = 16'h52b9; // 0x2a24
	13'h1513: q2 = 16'h0001; // 0x2a26
	13'h1514: q2 = 16'h75be; // 0x2a28
	13'h1515: q2 = 16'h4a9f; // 0x2a2a
	13'h1516: q2 = 16'h4cdf; // 0x2a2c
	13'h1517: q2 = 16'h00c0; // 0x2a2e
	13'h1518: q2 = 16'h4e5e; // 0x2a30
	13'h1519: q2 = 16'h4e75; // 0x2a32
	13'h151a: q2 = 16'h4e56; // 0x2a34
	13'h151b: q2 = 16'h0000; // 0x2a36
	13'h151c: q2 = 16'h48e7; // 0x2a38
	13'h151d: q2 = 16'h0304; // 0x2a3a
	13'h151e: q2 = 16'h2a7c; // 0x2a3c
	13'h151f: q2 = 16'h0001; // 0x2a3e
	13'h1520: q2 = 16'h759a; // 0x2a40
	13'h1521: q2 = 16'h4247; // 0x2a42
	13'h1522: q2 = 16'hbe7c; // 0x2a44
	13'h1523: q2 = 16'h000d; // 0x2a46
	13'h1524: q2 = 16'h6c08; // 0x2a48
	13'h1525: q2 = 16'h4295; // 0x2a4a
	13'h1526: q2 = 16'h5247; // 0x2a4c
	13'h1527: q2 = 16'h588d; // 0x2a4e
	13'h1528: q2 = 16'h60f2; // 0x2a50
	13'h1529: q2 = 16'h4a9f; // 0x2a52
	13'h152a: q2 = 16'h4cdf; // 0x2a54
	13'h152b: q2 = 16'h2080; // 0x2a56
	13'h152c: q2 = 16'h4e5e; // 0x2a58
	13'h152d: q2 = 16'h4e75; // 0x2a5a
	13'h152e: q2 = 16'h4e56; // 0x2a5c
	13'h152f: q2 = 16'hffdc; // 0x2a5e
	13'h1530: q2 = 16'h48e7; // 0x2a60
	13'h1531: q2 = 16'h3f00; // 0x2a62
	13'h1532: q2 = 16'h2639; // 0x2a64
	13'h1533: q2 = 16'h0001; // 0x2a66
	13'h1534: q2 = 16'h75ca; // 0x2a68
	13'h1535: q2 = 16'h4eb9; // 0x2a6a
	13'h1536: q2 = 16'h0000; // 0x2a6c
	13'h1537: q2 = 16'h0226; // 0x2a6e
	13'h1538: q2 = 16'h7e1f; // 0x2a70
	13'h1539: q2 = 16'hbe7c; // 0x2a72
	13'h153a: q2 = 16'h0004; // 0x2a74
	13'h153b: q2 = 16'h6d00; // 0x2a76
	13'h153c: q2 = 16'h02c4; // 0x2a78
	13'h153d: q2 = 16'h3ebc; // 0x2a7a
	13'h153e: q2 = 16'h001f; // 0x2a7c
	13'h153f: q2 = 16'h3007; // 0x2a7e
	13'h1540: q2 = 16'h9157; // 0x2a80
	13'h1541: q2 = 16'h0657; // 0x2a82
	13'h1542: q2 = 16'h003d; // 0x2a84
	13'h1543: q2 = 16'h200e; // 0x2a86
	13'h1544: q2 = 16'hd0bc; // 0x2a88
	13'h1545: q2 = 16'hffff; // 0x2a8a
	13'h1546: q2 = 16'hffdc; // 0x2a8c
	13'h1547: q2 = 16'h2f00; // 0x2a8e
	13'h1548: q2 = 16'h4eb9; // 0x2a90
	13'h1549: q2 = 16'h0000; // 0x2a92
	13'h154a: q2 = 16'h78f6; // 0x2a94
	13'h154b: q2 = 16'h4a9f; // 0x2a96
	13'h154c: q2 = 16'h0c2e; // 0x2a98
	13'h154d: q2 = 16'h0020; // 0x2a9a
	13'h154e: q2 = 16'hffdc; // 0x2a9c
	13'h154f: q2 = 16'h6604; // 0x2a9e
	13'h1550: q2 = 16'h7c02; // 0x2aa0
	13'h1551: q2 = 16'h6002; // 0x2aa2
	13'h1552: q2 = 16'h4246; // 0x2aa4
	13'h1553: q2 = 16'h701f; // 0x2aa6
	13'h1554: q2 = 16'h9047; // 0x2aa8
	13'h1555: q2 = 16'h48c0; // 0x2aaa
	13'h1556: q2 = 16'hd0bc; // 0x2aac
	13'h1557: q2 = 16'h0000; // 0x2aae
	13'h1558: q2 = 16'hfc5e; // 0x2ab0
	13'h1559: q2 = 16'h2040; // 0x2ab2
	13'h155a: q2 = 16'h1010; // 0x2ab4
	13'h155b: q2 = 16'h4880; // 0x2ab6
	13'h155c: q2 = 16'h3d40; // 0x2ab8
	13'h155d: q2 = 16'hfffe; // 0x2aba
	13'h155e: q2 = 16'h3eae; // 0x2abc
	13'h155f: q2 = 16'hfffe; // 0x2abe
	13'h1560: q2 = 16'h4267; // 0x2ac0
	13'h1561: q2 = 16'h3f06; // 0x2ac2
	13'h1562: q2 = 16'h3f07; // 0x2ac4
	13'h1563: q2 = 16'h200e; // 0x2ac6
	13'h1564: q2 = 16'hd0bc; // 0x2ac8
	13'h1565: q2 = 16'hffff; // 0x2aca
	13'h1566: q2 = 16'hffdc; // 0x2acc
	13'h1567: q2 = 16'h2f00; // 0x2ace
	13'h1568: q2 = 16'h4eb9; // 0x2ad0
	13'h1569: q2 = 16'h0000; // 0x2ad2
	13'h156a: q2 = 16'h026c; // 0x2ad4
	13'h156b: q2 = 16'hdefc; // 0x2ad6
	13'h156c: q2 = 16'h000a; // 0x2ad8
	13'h156d: q2 = 16'h7aff; // 0x2ada
	13'h156e: q2 = 16'h3007; // 0x2adc
	13'h156f: q2 = 16'h6000; // 0x2ade
	13'h1570: q2 = 16'h0198; // 0x2ae0
	13'h1571: q2 = 16'h2a39; // 0x2ae2
	13'h1572: q2 = 16'h0001; // 0x2ae4
	13'h1573: q2 = 16'h759a; // 0x2ae6
	13'h1574: q2 = 16'h6000; // 0x2ae8
	13'h1575: q2 = 16'h01a4; // 0x2aea
	13'h1576: q2 = 16'h2a39; // 0x2aec
	13'h1577: q2 = 16'h0001; // 0x2aee
	13'h1578: q2 = 16'h759e; // 0x2af0
	13'h1579: q2 = 16'h6000; // 0x2af2
	13'h157a: q2 = 16'h019a; // 0x2af4
	13'h157b: q2 = 16'h2f3c; // 0x2af6
	13'h157c: q2 = 16'h0000; // 0x2af8
	13'h157d: q2 = 16'h0002; // 0x2afa
	13'h157e: q2 = 16'h2f39; // 0x2afc
	13'h157f: q2 = 16'h0001; // 0x2afe
	13'h1580: q2 = 16'h759e; // 0x2b00
	13'h1581: q2 = 16'h4eb9; // 0x2b02
	13'h1582: q2 = 16'h0000; // 0x2b04
	13'h1583: q2 = 16'h7a50; // 0x2b06
	13'h1584: q2 = 16'hbf8f; // 0x2b08
	13'h1585: q2 = 16'h2a00; // 0x2b0a
	13'h1586: q2 = 16'hdab9; // 0x2b0c
	13'h1587: q2 = 16'h0001; // 0x2b0e
	13'h1588: q2 = 16'h759a; // 0x2b10
	13'h1589: q2 = 16'h6000; // 0x2b12
	13'h158a: q2 = 16'h017a; // 0x2b14
	13'h158b: q2 = 16'h2a39; // 0x2b16
	13'h158c: q2 = 16'h0001; // 0x2b18
	13'h158d: q2 = 16'h75a2; // 0x2b1a
	13'h158e: q2 = 16'h6000; // 0x2b1c
	13'h158f: q2 = 16'h0170; // 0x2b1e
	13'h1590: q2 = 16'h2a39; // 0x2b20
	13'h1591: q2 = 16'h0001; // 0x2b22
	13'h1592: q2 = 16'h75a6; // 0x2b24
	13'h1593: q2 = 16'h6000; // 0x2b26
	13'h1594: q2 = 16'h0166; // 0x2b28
	13'h1595: q2 = 16'h2a39; // 0x2b2a
	13'h1596: q2 = 16'h0001; // 0x2b2c
	13'h1597: q2 = 16'h75aa; // 0x2b2e
	13'h1598: q2 = 16'h6000; // 0x2b30
	13'h1599: q2 = 16'h015c; // 0x2b32
	13'h159a: q2 = 16'h2a39; // 0x2b34
	13'h159b: q2 = 16'h0001; // 0x2b36
	13'h159c: q2 = 16'h75ae; // 0x2b38
	13'h159d: q2 = 16'h6000; // 0x2b3a
	13'h159e: q2 = 16'h0152; // 0x2b3c
	13'h159f: q2 = 16'h2a39; // 0x2b3e
	13'h15a0: q2 = 16'h0001; // 0x2b40
	13'h15a1: q2 = 16'h75aa; // 0x2b42
	13'h15a2: q2 = 16'hdab9; // 0x2b44
	13'h15a3: q2 = 16'h0001; // 0x2b46
	13'h15a4: q2 = 16'h75ae; // 0x2b48
	13'h15a5: q2 = 16'h6000; // 0x2b4a
	13'h15a6: q2 = 16'h0142; // 0x2b4c
	13'h15a7: q2 = 16'h2a39; // 0x2b4e
	13'h15a8: q2 = 16'h0001; // 0x2b50
	13'h15a9: q2 = 16'h75b2; // 0x2b52
	13'h15aa: q2 = 16'h6000; // 0x2b54
	13'h15ab: q2 = 16'h0138; // 0x2b56
	13'h15ac: q2 = 16'h2a39; // 0x2b58
	13'h15ad: q2 = 16'h0001; // 0x2b5a
	13'h15ae: q2 = 16'h75b6; // 0x2b5c
	13'h15af: q2 = 16'h6000; // 0x2b5e
	13'h15b0: q2 = 16'h012e; // 0x2b60
	13'h15b1: q2 = 16'h2a39; // 0x2b62
	13'h15b2: q2 = 16'h0001; // 0x2b64
	13'h15b3: q2 = 16'h75ba; // 0x2b66
	13'h15b4: q2 = 16'h6000; // 0x2b68
	13'h15b5: q2 = 16'h0124; // 0x2b6a
	13'h15b6: q2 = 16'h2a39; // 0x2b6c
	13'h15b7: q2 = 16'h0001; // 0x2b6e
	13'h15b8: q2 = 16'h75b2; // 0x2b70
	13'h15b9: q2 = 16'hdab9; // 0x2b72
	13'h15ba: q2 = 16'h0001; // 0x2b74
	13'h15bb: q2 = 16'h75b6; // 0x2b76
	13'h15bc: q2 = 16'hdab9; // 0x2b78
	13'h15bd: q2 = 16'h0001; // 0x2b7a
	13'h15be: q2 = 16'h75ba; // 0x2b7c
	13'h15bf: q2 = 16'h6000; // 0x2b7e
	13'h15c0: q2 = 16'h010e; // 0x2b80
	13'h15c1: q2 = 16'h2f3c; // 0x2b82
	13'h15c2: q2 = 16'h0000; // 0x2b84
	13'h15c3: q2 = 16'h0002; // 0x2b86
	13'h15c4: q2 = 16'h2f39; // 0x2b88
	13'h15c5: q2 = 16'h0001; // 0x2b8a
	13'h15c6: q2 = 16'h759e; // 0x2b8c
	13'h15c7: q2 = 16'h4eb9; // 0x2b8e
	13'h15c8: q2 = 16'h0000; // 0x2b90
	13'h15c9: q2 = 16'h7a50; // 0x2b92
	13'h15ca: q2 = 16'hbf8f; // 0x2b94
	13'h15cb: q2 = 16'h2800; // 0x2b96
	13'h15cc: q2 = 16'hd8b9; // 0x2b98
	13'h15cd: q2 = 16'h0001; // 0x2b9a
	13'h15ce: q2 = 16'h759a; // 0x2b9c
	13'h15cf: q2 = 16'h4a84; // 0x2b9e
	13'h15d0: q2 = 16'h6604; // 0x2ba0
	13'h15d1: q2 = 16'h4285; // 0x2ba2
	13'h15d2: q2 = 16'h6024; // 0x2ba4
	13'h15d3: q2 = 16'h2f3c; // 0x2ba6
	13'h15d4: q2 = 16'h0000; // 0x2ba8
	13'h15d5: q2 = 16'h0064; // 0x2baa
	13'h15d6: q2 = 16'h2f39; // 0x2bac
	13'h15d7: q2 = 16'h0001; // 0x2bae
	13'h15d8: q2 = 16'h75be; // 0x2bb0
	13'h15d9: q2 = 16'h4eb9; // 0x2bb2
	13'h15da: q2 = 16'h0000; // 0x2bb4
	13'h15db: q2 = 16'h7a50; // 0x2bb6
	13'h15dc: q2 = 16'hbf8f; // 0x2bb8
	13'h15dd: q2 = 16'h2a00; // 0x2bba
	13'h15de: q2 = 16'h2f04; // 0x2bbc
	13'h15df: q2 = 16'h2f05; // 0x2bbe
	13'h15e0: q2 = 16'h4eb9; // 0x2bc0
	13'h15e1: q2 = 16'h0000; // 0x2bc2
	13'h15e2: q2 = 16'h79ac; // 0x2bc4
	13'h15e3: q2 = 16'hbf8f; // 0x2bc6
	13'h15e4: q2 = 16'h2a00; // 0x2bc8
	13'h15e5: q2 = 16'h6000; // 0x2bca
	13'h15e6: q2 = 16'h00c2; // 0x2bcc
	13'h15e7: q2 = 16'h2839; // 0x2bce
	13'h15e8: q2 = 16'h0001; // 0x2bd0
	13'h15e9: q2 = 16'h75aa; // 0x2bd2
	13'h15ea: q2 = 16'hd8b9; // 0x2bd4
	13'h15eb: q2 = 16'h0001; // 0x2bd6
	13'h15ec: q2 = 16'h75ae; // 0x2bd8
	13'h15ed: q2 = 16'h4a84; // 0x2bda
	13'h15ee: q2 = 16'h6604; // 0x2bdc
	13'h15ef: q2 = 16'h4285; // 0x2bde
	13'h15f0: q2 = 16'h600e; // 0x2be0
	13'h15f1: q2 = 16'h2f04; // 0x2be2
	13'h15f2: q2 = 16'h2f03; // 0x2be4
	13'h15f3: q2 = 16'h4eb9; // 0x2be6
	13'h15f4: q2 = 16'h0000; // 0x2be8
	13'h15f5: q2 = 16'h79ac; // 0x2bea
	13'h15f6: q2 = 16'hbf8f; // 0x2bec
	13'h15f7: q2 = 16'h2a00; // 0x2bee
	13'h15f8: q2 = 16'h6000; // 0x2bf0
	13'h15f9: q2 = 16'h009c; // 0x2bf2
	13'h15fa: q2 = 16'h2f3c; // 0x2bf4
	13'h15fb: q2 = 16'h0000; // 0x2bf6
	13'h15fc: q2 = 16'h0002; // 0x2bf8
	13'h15fd: q2 = 16'h2f39; // 0x2bfa
	13'h15fe: q2 = 16'h0001; // 0x2bfc
	13'h15ff: q2 = 16'h759e; // 0x2bfe
	13'h1600: q2 = 16'h4eb9; // 0x2c00
	13'h1601: q2 = 16'h0000; // 0x2c02
	13'h1602: q2 = 16'h7a50; // 0x2c04
	13'h1603: q2 = 16'hbf8f; // 0x2c06
	13'h1604: q2 = 16'h2800; // 0x2c08
	13'h1605: q2 = 16'hd8b9; // 0x2c0a
	13'h1606: q2 = 16'h0001; // 0x2c0c
	13'h1607: q2 = 16'h759a; // 0x2c0e
	13'h1608: q2 = 16'h4a84; // 0x2c10
	13'h1609: q2 = 16'h6604; // 0x2c12
	13'h160a: q2 = 16'h4285; // 0x2c14
	13'h160b: q2 = 16'h6012; // 0x2c16
	13'h160c: q2 = 16'h2f04; // 0x2c18
	13'h160d: q2 = 16'h2f39; // 0x2c1a
	13'h160e: q2 = 16'h0001; // 0x2c1c
	13'h160f: q2 = 16'h75c2; // 0x2c1e
	13'h1610: q2 = 16'h4eb9; // 0x2c20
	13'h1611: q2 = 16'h0000; // 0x2c22
	13'h1612: q2 = 16'h79ac; // 0x2c24
	13'h1613: q2 = 16'hbf8f; // 0x2c26
	13'h1614: q2 = 16'h2a00; // 0x2c28
	13'h1615: q2 = 16'h6062; // 0x2c2a
	13'h1616: q2 = 16'h2a39; // 0x2c2c
	13'h1617: q2 = 16'h0001; // 0x2c2e
	13'h1618: q2 = 16'h75c6; // 0x2c30
	13'h1619: q2 = 16'h605a; // 0x2c32
	13'h161a: q2 = 16'h2a03; // 0x2c34
	13'h161b: q2 = 16'h6056; // 0x2c36
	13'h161c: q2 = 16'h4a83; // 0x2c38
	13'h161d: q2 = 16'h6604; // 0x2c3a
	13'h161e: q2 = 16'h4285; // 0x2c3c
	13'h161f: q2 = 16'h6024; // 0x2c3e
	13'h1620: q2 = 16'h2f3c; // 0x2c40
	13'h1621: q2 = 16'h0000; // 0x2c42
	13'h1622: q2 = 16'h0064; // 0x2c44
	13'h1623: q2 = 16'h2f39; // 0x2c46
	13'h1624: q2 = 16'h0001; // 0x2c48
	13'h1625: q2 = 16'h75c2; // 0x2c4a
	13'h1626: q2 = 16'h4eb9; // 0x2c4c
	13'h1627: q2 = 16'h0000; // 0x2c4e
	13'h1628: q2 = 16'h7a50; // 0x2c50
	13'h1629: q2 = 16'hbf8f; // 0x2c52
	13'h162a: q2 = 16'h2a00; // 0x2c54
	13'h162b: q2 = 16'h2f03; // 0x2c56
	13'h162c: q2 = 16'h2f05; // 0x2c58
	13'h162d: q2 = 16'h4eb9; // 0x2c5a
	13'h162e: q2 = 16'h0000; // 0x2c5c
	13'h162f: q2 = 16'h79ac; // 0x2c5e
	13'h1630: q2 = 16'hbf8f; // 0x2c60
	13'h1631: q2 = 16'h2a00; // 0x2c62
	13'h1632: q2 = 16'h6028; // 0x2c64
	13'h1633: q2 = 16'h2a39; // 0x2c66
	13'h1634: q2 = 16'h0001; // 0x2c68
	13'h1635: q2 = 16'h75d2; // 0x2c6a
	13'h1636: q2 = 16'h6020; // 0x2c6c
	13'h1637: q2 = 16'h2a39; // 0x2c6e
	13'h1638: q2 = 16'h0001; // 0x2c70
	13'h1639: q2 = 16'h75ce; // 0x2c72
	13'h163a: q2 = 16'h6018; // 0x2c74
	13'h163b: q2 = 16'h6016; // 0x2c76
	13'h163c: q2 = 16'h5940; // 0x2c78
	13'h163d: q2 = 16'hb07c; // 0x2c7a
	13'h163e: q2 = 16'h0018; // 0x2c7c
	13'h163f: q2 = 16'h620e; // 0x2c7e
	13'h1640: q2 = 16'he540; // 0x2c80
	13'h1641: q2 = 16'h3040; // 0x2c82
	13'h1642: q2 = 16'hd1fc; // 0x2c84
	13'h1643: q2 = 16'h0000; // 0x2c86
	13'h1644: q2 = 16'hfc7a; // 0x2c88
	13'h1645: q2 = 16'h2050; // 0x2c8a
	13'h1646: q2 = 16'h4ed0; // 0x2c8c
	13'h1647: q2 = 16'hbabc; // 0x2c8e
	13'h1648: q2 = 16'hffff; // 0x2c90
	13'h1649: q2 = 16'hffff; // 0x2c92
	13'h164a: q2 = 16'h661a; // 0x2c94
	13'h164b: q2 = 16'h2ebc; // 0x2c96
	13'h164c: q2 = 16'h0000; // 0x2c98
	13'h164d: q2 = 16'hfcde; // 0x2c9a
	13'h164e: q2 = 16'h200e; // 0x2c9c
	13'h164f: q2 = 16'hd0bc; // 0x2c9e
	13'h1650: q2 = 16'hffff; // 0x2ca0
	13'h1651: q2 = 16'hffdc; // 0x2ca2
	13'h1652: q2 = 16'h2f00; // 0x2ca4
	13'h1653: q2 = 16'h4eb9; // 0x2ca6
	13'h1654: q2 = 16'h0000; // 0x2ca8
	13'h1655: q2 = 16'h0750; // 0x2caa
	13'h1656: q2 = 16'h4a9f; // 0x2cac
	13'h1657: q2 = 16'h603c; // 0x2cae
	13'h1658: q2 = 16'hbe7c; // 0x2cb0
	13'h1659: q2 = 16'h0007; // 0x2cb2
	13'h165a: q2 = 16'h6f06; // 0x2cb4
	13'h165b: q2 = 16'hbe7c; // 0x2cb6
	13'h165c: q2 = 16'h000d; // 0x2cb8
	13'h165d: q2 = 16'h6d06; // 0x2cba
	13'h165e: q2 = 16'hbe7c; // 0x2cbc
	13'h165f: q2 = 16'h0005; // 0x2cbe
	13'h1660: q2 = 16'h6616; // 0x2cc0
	13'h1661: q2 = 16'h200e; // 0x2cc2
	13'h1662: q2 = 16'hd0bc; // 0x2cc4
	13'h1663: q2 = 16'hffff; // 0x2cc6
	13'h1664: q2 = 16'hffdc; // 0x2cc8
	13'h1665: q2 = 16'h2e80; // 0x2cca
	13'h1666: q2 = 16'h2f05; // 0x2ccc
	13'h1667: q2 = 16'h4eb9; // 0x2cce
	13'h1668: q2 = 16'h0000; // 0x2cd0
	13'h1669: q2 = 16'hb976; // 0x2cd2
	13'h166a: q2 = 16'h4a9f; // 0x2cd4
	13'h166b: q2 = 16'h6014; // 0x2cd6
	13'h166c: q2 = 16'h200e; // 0x2cd8
	13'h166d: q2 = 16'hd0bc; // 0x2cda
	13'h166e: q2 = 16'hffff; // 0x2cdc
	13'h166f: q2 = 16'hffdc; // 0x2cde
	13'h1670: q2 = 16'h2e80; // 0x2ce0
	13'h1671: q2 = 16'h2f05; // 0x2ce2
	13'h1672: q2 = 16'h4eb9; // 0x2ce4
	13'h1673: q2 = 16'h0000; // 0x2ce6
	13'h1674: q2 = 16'h0892; // 0x2ce8
	13'h1675: q2 = 16'h4a9f; // 0x2cea
	13'h1676: q2 = 16'hbe7c; // 0x2cec
	13'h1677: q2 = 16'h000d; // 0x2cee
	13'h1678: q2 = 16'h6706; // 0x2cf0
	13'h1679: q2 = 16'hbe7c; // 0x2cf2
	13'h167a: q2 = 16'h0007; // 0x2cf4
	13'h167b: q2 = 16'h6618; // 0x2cf6
	13'h167c: q2 = 16'h2ebc; // 0x2cf8
	13'h167d: q2 = 16'h0000; // 0x2cfa
	13'h167e: q2 = 16'hfce0; // 0x2cfc
	13'h167f: q2 = 16'h200e; // 0x2cfe
	13'h1680: q2 = 16'hd0bc; // 0x2d00
	13'h1681: q2 = 16'hffff; // 0x2d02
	13'h1682: q2 = 16'hffdc; // 0x2d04
	13'h1683: q2 = 16'h2f00; // 0x2d06
	13'h1684: q2 = 16'h4eb9; // 0x2d08
	13'h1685: q2 = 16'h0000; // 0x2d0a
	13'h1686: q2 = 16'h0770; // 0x2d0c
	13'h1687: q2 = 16'h4a9f; // 0x2d0e
	13'h1688: q2 = 16'hbe7c; // 0x2d10
	13'h1689: q2 = 16'h001f; // 0x2d12
	13'h168a: q2 = 16'h6720; // 0x2d14
	13'h168b: q2 = 16'h3eae; // 0x2d16
	13'h168c: q2 = 16'hfffe; // 0x2d18
	13'h168d: q2 = 16'h4267; // 0x2d1a
	13'h168e: q2 = 16'h3f3c; // 0x2d1c
	13'h168f: q2 = 16'hffe1; // 0x2d1e
	13'h1690: q2 = 16'h3f07; // 0x2d20
	13'h1691: q2 = 16'h200e; // 0x2d22
	13'h1692: q2 = 16'hd0bc; // 0x2d24
	13'h1693: q2 = 16'hffff; // 0x2d26
	13'h1694: q2 = 16'hffdc; // 0x2d28
	13'h1695: q2 = 16'h2f00; // 0x2d2a
	13'h1696: q2 = 16'h4eb9; // 0x2d2c
	13'h1697: q2 = 16'h0000; // 0x2d2e
	13'h1698: q2 = 16'h026c; // 0x2d30
	13'h1699: q2 = 16'hdefc; // 0x2d32
	13'h169a: q2 = 16'h000a; // 0x2d34
	13'h169b: q2 = 16'h5347; // 0x2d36
	13'h169c: q2 = 16'h6000; // 0x2d38
	13'h169d: q2 = 16'hfd38; // 0x2d3a
	13'h169e: q2 = 16'h4a79; // 0x2d3c
	13'h169f: q2 = 16'h0001; // 0x2d3e
	13'h16a0: q2 = 16'h8a7e; // 0x2d40
	13'h16a1: q2 = 16'h6702; // 0x2d42
	13'h16a2: q2 = 16'h60f6; // 0x2d44
	13'h16a3: q2 = 16'h4a79; // 0x2d46
	13'h16a4: q2 = 16'h0001; // 0x2d48
	13'h16a5: q2 = 16'h8a7e; // 0x2d4a
	13'h16a6: q2 = 16'h6602; // 0x2d4c
	13'h16a7: q2 = 16'h60f6; // 0x2d4e
	13'h16a8: q2 = 16'h4a9f; // 0x2d50
	13'h16a9: q2 = 16'h4cdf; // 0x2d52
	13'h16aa: q2 = 16'h00f8; // 0x2d54
	13'h16ab: q2 = 16'h4e5e; // 0x2d56
	13'h16ac: q2 = 16'h4e75; // 0x2d58
	13'h16ad: q2 = 16'h4e56; // 0x2d5a
	13'h16ae: q2 = 16'h0000; // 0x2d5c
	13'h16af: q2 = 16'h48e7; // 0x2d5e
	13'h16b0: q2 = 16'h0300; // 0x2d60
	13'h16b1: q2 = 16'h2e39; // 0x2d62
	13'h16b2: q2 = 16'h0001; // 0x2d64
	13'h16b3: q2 = 16'h75ca; // 0x2d66
	13'h16b4: q2 = 16'h2007; // 0x2d68
	13'h16b5: q2 = 16'h90b9; // 0x2d6a
	13'h16b6: q2 = 16'h0001; // 0x2d6c
	13'h16b7: q2 = 16'h75d6; // 0x2d6e
	13'h16b8: q2 = 16'h7201; // 0x2d70
	13'h16b9: q2 = 16'h926e; // 0x2d72
	13'h16ba: q2 = 16'h0008; // 0x2d74
	13'h16bb: q2 = 16'he541; // 0x2d76
	13'h16bc: q2 = 16'h48c1; // 0x2d78
	13'h16bd: q2 = 16'hd2bc; // 0x2d7a
	13'h16be: q2 = 16'h0001; // 0x2d7c
	13'h16bf: q2 = 16'h75de; // 0x2d7e
	13'h16c0: q2 = 16'h2241; // 0x2d80
	13'h16c1: q2 = 16'hd191; // 0x2d82
	13'h16c2: q2 = 16'h23c7; // 0x2d84
	13'h16c3: q2 = 16'h0001; // 0x2d86
	13'h16c4: q2 = 16'h75d6; // 0x2d88
	13'h16c5: q2 = 16'h4a9f; // 0x2d8a
	13'h16c6: q2 = 16'h4cdf; // 0x2d8c
	13'h16c7: q2 = 16'h0080; // 0x2d8e
	13'h16c8: q2 = 16'h4e5e; // 0x2d90
	13'h16c9: q2 = 16'h4e75; // 0x2d92
	13'h16ca: q2 = 16'h4e56; // 0x2d94
	13'h16cb: q2 = 16'hff2c; // 0x2d96
	13'h16cc: q2 = 16'h48e7; // 0x2d98
	13'h16cd: q2 = 16'h1f1c; // 0x2d9a
	13'h16ce: q2 = 16'h7001; // 0x2d9c
	13'h16cf: q2 = 16'h9079; // 0x2d9e
	13'h16d0: q2 = 16'h0001; // 0x2da0
	13'h16d1: q2 = 16'h805a; // 0x2da2
	13'h16d2: q2 = 16'h33c0; // 0x2da4
	13'h16d3: q2 = 16'h0001; // 0x2da6
	13'h16d4: q2 = 16'h805a; // 0x2da8
	13'h16d5: q2 = 16'h4a79; // 0x2daa
	13'h16d6: q2 = 16'h0001; // 0x2dac
	13'h16d7: q2 = 16'h805a; // 0x2dae
	13'h16d8: q2 = 16'h6700; // 0x2db0
	13'h16d9: q2 = 16'h04f2; // 0x2db2
	13'h16da: q2 = 16'h4246; // 0x2db4
	13'h16db: q2 = 16'h287c; // 0x2db6
	13'h16dc: q2 = 16'h0001; // 0x2db8
	13'h16dd: q2 = 16'h8072; // 0x2dba
	13'h16de: q2 = 16'hbc7c; // 0x2dbc
	13'h16df: q2 = 16'h0030; // 0x2dbe
	13'h16e0: q2 = 16'h6c0c; // 0x2dc0
	13'h16e1: q2 = 16'h026c; // 0x2dc2
	13'h16e2: q2 = 16'h00df; // 0x2dc4
	13'h16e3: q2 = 16'h0006; // 0x2dc6
	13'h16e4: q2 = 16'h5246; // 0x2dc8
	13'h16e5: q2 = 16'h508c; // 0x2dca
	13'h16e6: q2 = 16'h60ee; // 0x2dcc
	13'h16e7: q2 = 16'h4246; // 0x2dce
	13'h16e8: q2 = 16'h2d7c; // 0x2dd0
	13'h16e9: q2 = 16'h0001; // 0x2dd2
	13'h16ea: q2 = 16'h893e; // 0x2dd4
	13'h16eb: q2 = 16'hfffc; // 0x2dd6
	13'h16ec: q2 = 16'hbc79; // 0x2dd8
	13'h16ed: q2 = 16'h0001; // 0x2dda
	13'h16ee: q2 = 16'h7fa8; // 0x2ddc
	13'h16ef: q2 = 16'h6c00; // 0x2dde
	13'h16f0: q2 = 16'h00d6; // 0x2de0
	13'h16f1: q2 = 16'h287c; // 0x2de2
	13'h16f2: q2 = 16'h0001; // 0x2de4
	13'h16f3: q2 = 16'h8072; // 0x2de6
	13'h16f4: q2 = 16'h3014; // 0x2de8
	13'h16f5: q2 = 16'h226e; // 0x2dea
	13'h16f6: q2 = 16'hfffc; // 0x2dec
	13'h16f7: q2 = 16'h9051; // 0x2dee
	13'h16f8: q2 = 16'h3e00; // 0x2df0
	13'h16f9: q2 = 16'h4a47; // 0x2df2
	13'h16fa: q2 = 16'h6c06; // 0x2df4
	13'h16fb: q2 = 16'h3007; // 0x2df6
	13'h16fc: q2 = 16'h4440; // 0x2df8
	13'h16fd: q2 = 16'h3e00; // 0x2dfa
	13'h16fe: q2 = 16'hbe7c; // 0x2dfc
	13'h16ff: q2 = 16'h0800; // 0x2dfe
	13'h1700: q2 = 16'h6c22; // 0x2e00
	13'h1701: q2 = 16'h302c; // 0x2e02
	13'h1702: q2 = 16'h0002; // 0x2e04
	13'h1703: q2 = 16'h226e; // 0x2e06
	13'h1704: q2 = 16'hfffc; // 0x2e08
	13'h1705: q2 = 16'h9069; // 0x2e0a
	13'h1706: q2 = 16'h0002; // 0x2e0c
	13'h1707: q2 = 16'h3e00; // 0x2e0e
	13'h1708: q2 = 16'h9e7c; // 0x2e10
	13'h1709: q2 = 16'h0080; // 0x2e12
	13'h170a: q2 = 16'h4a47; // 0x2e14
	13'h170b: q2 = 16'h6f0c; // 0x2e16
	13'h170c: q2 = 16'hbe7c; // 0x2e18
	13'h170d: q2 = 16'h0800; // 0x2e1a
	13'h170e: q2 = 16'h6c06; // 0x2e1c
	13'h170f: q2 = 16'h006c; // 0x2e1e
	13'h1710: q2 = 16'h0020; // 0x2e20
	13'h1711: q2 = 16'h0006; // 0x2e22
	13'h1712: q2 = 16'h082c; // 0x2e24
	13'h1713: q2 = 16'h0005; // 0x2e26
	13'h1714: q2 = 16'h0007; // 0x2e28
	13'h1715: q2 = 16'h6700; // 0x2e2a
	13'h1716: q2 = 16'h007c; // 0x2e2c
	13'h1717: q2 = 16'h206e; // 0x2e2e
	13'h1718: q2 = 16'hfffc; // 0x2e30
	13'h1719: q2 = 16'h3028; // 0x2e32
	13'h171a: q2 = 16'h0002; // 0x2e34
	13'h171b: q2 = 16'hd07c; // 0x2e36
	13'h171c: q2 = 16'h0380; // 0x2e38
	13'h171d: q2 = 16'hb06c; // 0x2e3a
	13'h171e: q2 = 16'h0002; // 0x2e3c
	13'h171f: q2 = 16'h6f10; // 0x2e3e
	13'h1720: q2 = 16'h0079; // 0x2e40
	13'h1721: q2 = 16'h0020; // 0x2e42
	13'h1722: q2 = 16'h0001; // 0x2e44
	13'h1723: q2 = 16'h8080; // 0x2e46
	13'h1724: q2 = 16'h0079; // 0x2e48
	13'h1725: q2 = 16'h0020; // 0x2e4a
	13'h1726: q2 = 16'h0001; // 0x2e4c
	13'h1727: q2 = 16'h80a8; // 0x2e4e
	13'h1728: q2 = 16'h4ab9; // 0x2e50
	13'h1729: q2 = 16'h0001; // 0x2e52
	13'h172a: q2 = 16'h7f36; // 0x2e54
	13'h172b: q2 = 16'h672e; // 0x2e56
	13'h172c: q2 = 16'h2079; // 0x2e58
	13'h172d: q2 = 16'h0001; // 0x2e5a
	13'h172e: q2 = 16'h7f36; // 0x2e5c
	13'h172f: q2 = 16'h2068; // 0x2e5e
	13'h1730: q2 = 16'h0012; // 0x2e60
	13'h1731: q2 = 16'h3028; // 0x2e62
	13'h1732: q2 = 16'h0002; // 0x2e64
	13'h1733: q2 = 16'h226e; // 0x2e66
	13'h1734: q2 = 16'hfffc; // 0x2e68
	13'h1735: q2 = 16'h3229; // 0x2e6a
	13'h1736: q2 = 16'h0002; // 0x2e6c
	13'h1737: q2 = 16'hd27c; // 0x2e6e
	13'h1738: q2 = 16'h0380; // 0x2e70
	13'h1739: q2 = 16'hb041; // 0x2e72
	13'h173a: q2 = 16'h6c10; // 0x2e74
	13'h173b: q2 = 16'h7020; // 0x2e76
	13'h173c: q2 = 16'h2279; // 0x2e78
	13'h173d: q2 = 16'h0001; // 0x2e7a
	13'h173e: q2 = 16'h7f36; // 0x2e7c
	13'h173f: q2 = 16'h2269; // 0x2e7e
	13'h1740: q2 = 16'h0012; // 0x2e80
	13'h1741: q2 = 16'h8169; // 0x2e82
	13'h1742: q2 = 16'h0006; // 0x2e84
	13'h1743: q2 = 16'h4ab9; // 0x2e86
	13'h1744: q2 = 16'h0001; // 0x2e88
	13'h1745: q2 = 16'h7f32; // 0x2e8a
	13'h1746: q2 = 16'h6710; // 0x2e8c
	13'h1747: q2 = 16'h7020; // 0x2e8e
	13'h1748: q2 = 16'h2279; // 0x2e90
	13'h1749: q2 = 16'h0001; // 0x2e92
	13'h174a: q2 = 16'h7f32; // 0x2e94
	13'h174b: q2 = 16'h2269; // 0x2e96
	13'h174c: q2 = 16'h0012; // 0x2e98
	13'h174d: q2 = 16'h8169; // 0x2e9a
	13'h174e: q2 = 16'h0006; // 0x2e9c
	13'h174f: q2 = 16'h0079; // 0x2e9e
	13'h1750: q2 = 16'h0020; // 0x2ea0
	13'h1751: q2 = 16'h0001; // 0x2ea2
	13'h1752: q2 = 16'h80a0; // 0x2ea4
	13'h1753: q2 = 16'h600e; // 0x2ea6
	13'h1754: q2 = 16'h5246; // 0x2ea8
	13'h1755: q2 = 16'h06ae; // 0x2eaa
	13'h1756: q2 = 16'h0000; // 0x2eac
	13'h1757: q2 = 16'h0010; // 0x2eae
	13'h1758: q2 = 16'hfffc; // 0x2eb0
	13'h1759: q2 = 16'h6000; // 0x2eb2
	13'h175a: q2 = 16'hff24; // 0x2eb4
	13'h175b: q2 = 16'h7a08; // 0x2eb6
	13'h175c: q2 = 16'h2d7c; // 0x2eb8
	13'h175d: q2 = 16'h0001; // 0x2eba
	13'h175e: q2 = 16'h89be; // 0x2ebc
	13'h175f: q2 = 16'hfff8; // 0x2ebe
	13'h1760: q2 = 16'h287c; // 0x2ec0
	13'h1761: q2 = 16'h0001; // 0x2ec2
	13'h1762: q2 = 16'h80b2; // 0x2ec4
	13'h1763: q2 = 16'hba7c; // 0x2ec6
	13'h1764: q2 = 16'h000b; // 0x2ec8
	13'h1765: q2 = 16'h6e00; // 0x2eca
	13'h1766: q2 = 16'h00b2; // 0x2ecc
	13'h1767: q2 = 16'h206e; // 0x2ece
	13'h1768: q2 = 16'hfff8; // 0x2ed0
	13'h1769: q2 = 16'h3828; // 0x2ed2
	13'h176a: q2 = 16'h0018; // 0x2ed4
	13'h176b: q2 = 16'h4246; // 0x2ed6
	13'h176c: q2 = 16'h2d7c; // 0x2ed8
	13'h176d: q2 = 16'h0001; // 0x2eda
	13'h176e: q2 = 16'h893e; // 0x2edc
	13'h176f: q2 = 16'hfffc; // 0x2ede
	13'h1770: q2 = 16'hbc79; // 0x2ee0
	13'h1771: q2 = 16'h0001; // 0x2ee2
	13'h1772: q2 = 16'h7fa8; // 0x2ee4
	13'h1773: q2 = 16'h6c00; // 0x2ee6
	13'h1774: q2 = 16'h0086; // 0x2ee8
	13'h1775: q2 = 16'h3014; // 0x2eea
	13'h1776: q2 = 16'h226e; // 0x2eec
	13'h1777: q2 = 16'hfffc; // 0x2eee
	13'h1778: q2 = 16'h9051; // 0x2ef0
	13'h1779: q2 = 16'h3e00; // 0x2ef2
	13'h177a: q2 = 16'h4a47; // 0x2ef4
	13'h177b: q2 = 16'h6c06; // 0x2ef6
	13'h177c: q2 = 16'h3007; // 0x2ef8
	13'h177d: q2 = 16'h4440; // 0x2efa
	13'h177e: q2 = 16'h3e00; // 0x2efc
	13'h177f: q2 = 16'hbe7c; // 0x2efe
	13'h1780: q2 = 16'h0800; // 0x2f00
	13'h1781: q2 = 16'h6c5c; // 0x2f02
	13'h1782: q2 = 16'h3004; // 0x2f04
	13'h1783: q2 = 16'h226e; // 0x2f06
	13'h1784: q2 = 16'hfffc; // 0x2f08
	13'h1785: q2 = 16'h9069; // 0x2f0a
	13'h1786: q2 = 16'h0002; // 0x2f0c
	13'h1787: q2 = 16'h3e00; // 0x2f0e
	13'h1788: q2 = 16'hde7c; // 0x2f10
	13'h1789: q2 = 16'hff80; // 0x2f12
	13'h178a: q2 = 16'h4a47; // 0x2f14
	13'h178b: q2 = 16'h6f48; // 0x2f16
	13'h178c: q2 = 16'hbe7c; // 0x2f18
	13'h178d: q2 = 16'h0800; // 0x2f1a
	13'h178e: q2 = 16'h6c42; // 0x2f1c
	13'h178f: q2 = 16'h006c; // 0x2f1e
	13'h1790: q2 = 16'h0020; // 0x2f20
	13'h1791: q2 = 16'h0006; // 0x2f22
	13'h1792: q2 = 16'h006c; // 0x2f24
	13'h1793: q2 = 16'h0020; // 0x2f26
	13'h1794: q2 = 16'h0026; // 0x2f28
	13'h1795: q2 = 16'h206e; // 0x2f2a
	13'h1796: q2 = 16'hfffc; // 0x2f2c
	13'h1797: q2 = 16'h3028; // 0x2f2e
	13'h1798: q2 = 16'h0002; // 0x2f30
	13'h1799: q2 = 16'hd07c; // 0x2f32
	13'h179a: q2 = 16'h0380; // 0x2f34
	13'h179b: q2 = 16'hb06c; // 0x2f36
	13'h179c: q2 = 16'h0002; // 0x2f38
	13'h179d: q2 = 16'h6f06; // 0x2f3a
	13'h179e: q2 = 16'h006c; // 0x2f3c
	13'h179f: q2 = 16'h0020; // 0x2f3e
	13'h17a0: q2 = 16'h0046; // 0x2f40
	13'h17a1: q2 = 16'h206e; // 0x2f42
	13'h17a2: q2 = 16'hfff8; // 0x2f44
	13'h17a3: q2 = 16'h4aa8; // 0x2f46
	13'h17a4: q2 = 16'h0010; // 0x2f48
	13'h17a5: q2 = 16'h6712; // 0x2f4a
	13'h17a6: q2 = 16'h7020; // 0x2f4c
	13'h17a7: q2 = 16'h226e; // 0x2f4e
	13'h17a8: q2 = 16'hfff8; // 0x2f50
	13'h17a9: q2 = 16'h2269; // 0x2f52
	13'h17aa: q2 = 16'h0010; // 0x2f54
	13'h17ab: q2 = 16'h2269; // 0x2f56
	13'h17ac: q2 = 16'h0012; // 0x2f58
	13'h17ad: q2 = 16'h8169; // 0x2f5a
	13'h17ae: q2 = 16'h0006; // 0x2f5c
	13'h17af: q2 = 16'h600e; // 0x2f5e
	13'h17b0: q2 = 16'h5246; // 0x2f60
	13'h17b1: q2 = 16'h06ae; // 0x2f62
	13'h17b2: q2 = 16'h0000; // 0x2f64
	13'h17b3: q2 = 16'h0010; // 0x2f66
	13'h17b4: q2 = 16'hfffc; // 0x2f68
	13'h17b5: q2 = 16'h6000; // 0x2f6a
	13'h17b6: q2 = 16'hff74; // 0x2f6c
	13'h17b7: q2 = 16'h5245; // 0x2f6e
	13'h17b8: q2 = 16'h06ae; // 0x2f70
	13'h17b9: q2 = 16'h0000; // 0x2f72
	13'h17ba: q2 = 16'h002e; // 0x2f74
	13'h17bb: q2 = 16'hfff8; // 0x2f76
	13'h17bc: q2 = 16'h508c; // 0x2f78
	13'h17bd: q2 = 16'h6000; // 0x2f7a
	13'h17be: q2 = 16'hff4a; // 0x2f7c
	13'h17bf: q2 = 16'h4a79; // 0x2f7e
	13'h17c0: q2 = 16'h0001; // 0x2f80
	13'h17c1: q2 = 16'h7faa; // 0x2f82
	13'h17c2: q2 = 16'h6742; // 0x2f84
	13'h17c3: q2 = 16'h7a14; // 0x2f86
	13'h17c4: q2 = 16'h2d7c; // 0x2f88
	13'h17c5: q2 = 16'h0001; // 0x2f8a
	13'h17c6: q2 = 16'h7bda; // 0x2f8c
	13'h17c7: q2 = 16'hfff0; // 0x2f8e
	13'h17c8: q2 = 16'h287c; // 0x2f90
	13'h17c9: q2 = 16'h0001; // 0x2f92
	13'h17ca: q2 = 16'h8112; // 0x2f94
	13'h17cb: q2 = 16'hba7c; // 0x2f96
	13'h17cc: q2 = 16'h002d; // 0x2f98
	13'h17cd: q2 = 16'h6e2c; // 0x2f9a
	13'h17ce: q2 = 16'h206e; // 0x2f9c
	13'h17cf: q2 = 16'hfff0; // 0x2f9e
	13'h17d0: q2 = 16'h0c68; // 0x2fa0
	13'h17d1: q2 = 16'h0006; // 0x2fa2
	13'h17d2: q2 = 16'h0008; // 0x2fa4
	13'h17d3: q2 = 16'h6612; // 0x2fa6
	13'h17d4: q2 = 16'h206e; // 0x2fa8
	13'h17d5: q2 = 16'hfff0; // 0x2faa
	13'h17d6: q2 = 16'h0c68; // 0x2fac
	13'h17d7: q2 = 16'h0001; // 0x2fae
	13'h17d8: q2 = 16'h001a; // 0x2fb0
	13'h17d9: q2 = 16'h6606; // 0x2fb2
	13'h17da: q2 = 16'h006c; // 0x2fb4
	13'h17db: q2 = 16'h0020; // 0x2fb6
	13'h17dc: q2 = 16'h0006; // 0x2fb8
	13'h17dd: q2 = 16'h5245; // 0x2fba
	13'h17de: q2 = 16'h06ae; // 0x2fbc
	13'h17df: q2 = 16'h0000; // 0x2fbe
	13'h17e0: q2 = 16'h001c; // 0x2fc0
	13'h17e1: q2 = 16'hfff0; // 0x2fc2
	13'h17e2: q2 = 16'h508c; // 0x2fc4
	13'h17e3: q2 = 16'h60ce; // 0x2fc6
	13'h17e4: q2 = 16'h47ee; // 0x2fc8
	13'h17e5: q2 = 16'hff2c; // 0x2fca
	13'h17e6: q2 = 16'h4246; // 0x2fcc
	13'h17e7: q2 = 16'h41ee; // 0x2fce
	13'h17e8: q2 = 16'hff90; // 0x2fd0
	13'h17e9: q2 = 16'h2d48; // 0x2fd2
	13'h17ea: q2 = 16'hff8c; // 0x2fd4
	13'h17eb: q2 = 16'hbc7c; // 0x2fd6
	13'h17ec: q2 = 16'h0030; // 0x2fd8
	13'h17ed: q2 = 16'h6c0e; // 0x2fda
	13'h17ee: q2 = 16'h206e; // 0x2fdc
	13'h17ef: q2 = 16'hff8c; // 0x2fde
	13'h17f0: q2 = 16'h4250; // 0x2fe0
	13'h17f1: q2 = 16'h5246; // 0x2fe2
	13'h17f2: q2 = 16'h54ae; // 0x2fe4
	13'h17f3: q2 = 16'hff8c; // 0x2fe6
	13'h17f4: q2 = 16'h60ec; // 0x2fe8
	13'h17f5: q2 = 16'h7aff; // 0x2fea
	13'h17f6: q2 = 16'h3039; // 0x2fec
	13'h17f7: q2 = 16'h0001; // 0x2fee
	13'h17f8: q2 = 16'h8074; // 0x2ff0
	13'h17f9: q2 = 16'hb045; // 0x2ff2
	13'h17fa: q2 = 16'h6d0e; // 0x2ff4
	13'h17fb: q2 = 16'h4a6e; // 0x2ff6
	13'h17fc: q2 = 16'hff90; // 0x2ff8
	13'h17fd: q2 = 16'h6608; // 0x2ffa
	13'h17fe: q2 = 16'h3a39; // 0x2ffc
	13'h17ff: q2 = 16'h0001; // 0x2ffe
	13'h1800: q2 = 16'h8074; // 0x3000
	13'h1801: q2 = 16'h4247; // 0x3002
	13'h1802: q2 = 16'h7c08; // 0x3004
	13'h1803: q2 = 16'h2d7c; // 0x3006
	13'h1804: q2 = 16'h0001; // 0x3008
	13'h1805: q2 = 16'h89be; // 0x300a
	13'h1806: q2 = 16'hfff8; // 0x300c
	13'h1807: q2 = 16'hbc7c; // 0x300e
	13'h1808: q2 = 16'h000b; // 0x3010
	13'h1809: q2 = 16'h6e32; // 0x3012
	13'h180a: q2 = 16'h206e; // 0x3014
	13'h180b: q2 = 16'hfff8; // 0x3016
	13'h180c: q2 = 16'h3828; // 0x3018
	13'h180d: q2 = 16'h0018; // 0x301a
	13'h180e: q2 = 16'hb845; // 0x301c
	13'h180f: q2 = 16'h6d1a; // 0x301e
	13'h1810: q2 = 16'h3006; // 0x3020
	13'h1811: q2 = 16'he340; // 0x3022
	13'h1812: q2 = 16'h48c0; // 0x3024
	13'h1813: q2 = 16'hd08e; // 0x3026
	13'h1814: q2 = 16'h2040; // 0x3028
	13'h1815: q2 = 16'h4a68; // 0x302a
	13'h1816: q2 = 16'hff90; // 0x302c
	13'h1817: q2 = 16'h660a; // 0x302e
	13'h1818: q2 = 16'h3a04; // 0x3030
	13'h1819: q2 = 16'h3e06; // 0x3032
	13'h181a: q2 = 16'h2d6e; // 0x3034
	13'h181b: q2 = 16'hfff8; // 0x3036
	13'h181c: q2 = 16'hfff4; // 0x3038
	13'h181d: q2 = 16'h5246; // 0x303a
	13'h181e: q2 = 16'h06ae; // 0x303c
	13'h181f: q2 = 16'h0000; // 0x303e
	13'h1820: q2 = 16'h002e; // 0x3040
	13'h1821: q2 = 16'hfff8; // 0x3042
	13'h1822: q2 = 16'h60c8; // 0x3044
	13'h1823: q2 = 16'hba7c; // 0x3046
	13'h1824: q2 = 16'hffff; // 0x3048
	13'h1825: q2 = 16'h6700; // 0x304a
	13'h1826: q2 = 16'h0166; // 0x304c
	13'h1827: q2 = 16'h4a47; // 0x304e
	13'h1828: q2 = 16'h6600; // 0x3050
	13'h1829: q2 = 16'h00d6; // 0x3052
	13'h182a: q2 = 16'h3687; // 0x3054
	13'h182b: q2 = 16'h548b; // 0x3056
	13'h182c: q2 = 16'h3007; // 0x3058
	13'h182d: q2 = 16'he340; // 0x305a
	13'h182e: q2 = 16'h48c0; // 0x305c
	13'h182f: q2 = 16'hd08e; // 0x305e
	13'h1830: q2 = 16'h2040; // 0x3060
	13'h1831: q2 = 16'h317c; // 0x3062
	13'h1832: q2 = 16'h0001; // 0x3064
	13'h1833: q2 = 16'hff90; // 0x3066
	13'h1834: q2 = 16'h7c01; // 0x3068
	13'h1835: q2 = 16'hbc7c; // 0x306a
	13'h1836: q2 = 16'h0004; // 0x306c
	13'h1837: q2 = 16'h6e18; // 0x306e
	13'h1838: q2 = 16'h3686; // 0x3070
	13'h1839: q2 = 16'h548b; // 0x3072
	13'h183a: q2 = 16'h3006; // 0x3074
	13'h183b: q2 = 16'he340; // 0x3076
	13'h183c: q2 = 16'h48c0; // 0x3078
	13'h183d: q2 = 16'hd08e; // 0x307a
	13'h183e: q2 = 16'h2040; // 0x307c
	13'h183f: q2 = 16'h317c; // 0x307e
	13'h1840: q2 = 16'h0001; // 0x3080
	13'h1841: q2 = 16'hff90; // 0x3082
	13'h1842: q2 = 16'h5246; // 0x3084
	13'h1843: q2 = 16'h60e2; // 0x3086
	13'h1844: q2 = 16'h36bc; // 0x3088
	13'h1845: q2 = 16'h0006; // 0x308a
	13'h1846: q2 = 16'h548b; // 0x308c
	13'h1847: q2 = 16'h3d7c; // 0x308e
	13'h1848: q2 = 16'h0001; // 0x3090
	13'h1849: q2 = 16'hff9c; // 0x3092
	13'h184a: q2 = 16'h36bc; // 0x3094
	13'h184b: q2 = 16'h0005; // 0x3096
	13'h184c: q2 = 16'h548b; // 0x3098
	13'h184d: q2 = 16'h3d7c; // 0x309a
	13'h184e: q2 = 16'h0001; // 0x309c
	13'h184f: q2 = 16'hff9a; // 0x309e
	13'h1850: q2 = 16'h36bc; // 0x30a0
	13'h1851: q2 = 16'h0007; // 0x30a2
	13'h1852: q2 = 16'h548b; // 0x30a4
	13'h1853: q2 = 16'h3d7c; // 0x30a6
	13'h1854: q2 = 16'h0001; // 0x30a8
	13'h1855: q2 = 16'hff9e; // 0x30aa
	13'h1856: q2 = 16'h4ab9; // 0x30ac
	13'h1857: q2 = 16'h0001; // 0x30ae
	13'h1858: q2 = 16'h7f32; // 0x30b0
	13'h1859: q2 = 16'h6734; // 0x30b2
	13'h185a: q2 = 16'h2079; // 0x30b4
	13'h185b: q2 = 16'h0001; // 0x30b6
	13'h185c: q2 = 16'h7f32; // 0x30b8
	13'h185d: q2 = 16'h2028; // 0x30ba
	13'h185e: q2 = 16'h0012; // 0x30bc
	13'h185f: q2 = 16'h90bc; // 0x30be
	13'h1860: q2 = 16'h0001; // 0x30c0
	13'h1861: q2 = 16'h8072; // 0x30c2
	13'h1862: q2 = 16'he680; // 0x30c4
	13'h1863: q2 = 16'h3680; // 0x30c6
	13'h1864: q2 = 16'h548b; // 0x30c8
	13'h1865: q2 = 16'h2079; // 0x30ca
	13'h1866: q2 = 16'h0001; // 0x30cc
	13'h1867: q2 = 16'h7f32; // 0x30ce
	13'h1868: q2 = 16'h2028; // 0x30d0
	13'h1869: q2 = 16'h0012; // 0x30d2
	13'h186a: q2 = 16'h90bc; // 0x30d4
	13'h186b: q2 = 16'h0001; // 0x30d6
	13'h186c: q2 = 16'h8072; // 0x30d8
	13'h186d: q2 = 16'he680; // 0x30da
	13'h186e: q2 = 16'he380; // 0x30dc
	13'h186f: q2 = 16'hd08e; // 0x30de
	13'h1870: q2 = 16'h2040; // 0x30e0
	13'h1871: q2 = 16'h317c; // 0x30e2
	13'h1872: q2 = 16'h0001; // 0x30e4
	13'h1873: q2 = 16'hff90; // 0x30e6
	13'h1874: q2 = 16'h4ab9; // 0x30e8
	13'h1875: q2 = 16'h0001; // 0x30ea
	13'h1876: q2 = 16'h7f36; // 0x30ec
	13'h1877: q2 = 16'h6734; // 0x30ee
	13'h1878: q2 = 16'h2079; // 0x30f0
	13'h1879: q2 = 16'h0001; // 0x30f2
	13'h187a: q2 = 16'h7f36; // 0x30f4
	13'h187b: q2 = 16'h2028; // 0x30f6
	13'h187c: q2 = 16'h0012; // 0x30f8
	13'h187d: q2 = 16'h90bc; // 0x30fa
	13'h187e: q2 = 16'h0001; // 0x30fc
	13'h187f: q2 = 16'h8072; // 0x30fe
	13'h1880: q2 = 16'he680; // 0x3100
	13'h1881: q2 = 16'h3680; // 0x3102
	13'h1882: q2 = 16'h548b; // 0x3104
	13'h1883: q2 = 16'h2079; // 0x3106
	13'h1884: q2 = 16'h0001; // 0x3108
	13'h1885: q2 = 16'h7f36; // 0x310a
	13'h1886: q2 = 16'h2028; // 0x310c
	13'h1887: q2 = 16'h0012; // 0x310e
	13'h1888: q2 = 16'h90bc; // 0x3110
	13'h1889: q2 = 16'h0001; // 0x3112
	13'h188a: q2 = 16'h8072; // 0x3114
	13'h188b: q2 = 16'he680; // 0x3116
	13'h188c: q2 = 16'he380; // 0x3118
	13'h188d: q2 = 16'hd08e; // 0x311a
	13'h188e: q2 = 16'h2040; // 0x311c
	13'h188f: q2 = 16'h317c; // 0x311e
	13'h1890: q2 = 16'h0001; // 0x3120
	13'h1891: q2 = 16'hff90; // 0x3122
	13'h1892: q2 = 16'h6000; // 0x3124
	13'h1893: q2 = 16'h0088; // 0x3126
	13'h1894: q2 = 16'h3687; // 0x3128
	13'h1895: q2 = 16'h548b; // 0x312a
	13'h1896: q2 = 16'h3007; // 0x312c
	13'h1897: q2 = 16'he340; // 0x312e
	13'h1898: q2 = 16'h48c0; // 0x3130
	13'h1899: q2 = 16'hd08e; // 0x3132
	13'h189a: q2 = 16'h2040; // 0x3134
	13'h189b: q2 = 16'h317c; // 0x3136
	13'h189c: q2 = 16'h0001; // 0x3138
	13'h189d: q2 = 16'hff90; // 0x313a
	13'h189e: q2 = 16'h3007; // 0x313c
	13'h189f: q2 = 16'h5840; // 0x313e
	13'h18a0: q2 = 16'h3680; // 0x3140
	13'h18a1: q2 = 16'h548b; // 0x3142
	13'h18a2: q2 = 16'h3007; // 0x3144
	13'h18a3: q2 = 16'he340; // 0x3146
	13'h18a4: q2 = 16'h48c0; // 0x3148
	13'h18a5: q2 = 16'hd08e; // 0x314a
	13'h18a6: q2 = 16'h2040; // 0x314c
	13'h18a7: q2 = 16'h317c; // 0x314e
	13'h18a8: q2 = 16'h0001; // 0x3150
	13'h18a9: q2 = 16'hff98; // 0x3152
	13'h18aa: q2 = 16'h3007; // 0x3154
	13'h18ab: q2 = 16'h5040; // 0x3156
	13'h18ac: q2 = 16'h3680; // 0x3158
	13'h18ad: q2 = 16'h548b; // 0x315a
	13'h18ae: q2 = 16'h3007; // 0x315c
	13'h18af: q2 = 16'he340; // 0x315e
	13'h18b0: q2 = 16'h48c0; // 0x3160
	13'h18b1: q2 = 16'hd08e; // 0x3162
	13'h18b2: q2 = 16'h2040; // 0x3164
	13'h18b3: q2 = 16'h317c; // 0x3166
	13'h18b4: q2 = 16'h0001; // 0x3168
	13'h18b5: q2 = 16'hffa0; // 0x316a
	13'h18b6: q2 = 16'h206e; // 0x316c
	13'h18b7: q2 = 16'hfff4; // 0x316e
	13'h18b8: q2 = 16'h4aa8; // 0x3170
	13'h18b9: q2 = 16'h0010; // 0x3172
	13'h18ba: q2 = 16'h6738; // 0x3174
	13'h18bb: q2 = 16'h206e; // 0x3176
	13'h18bc: q2 = 16'hfff4; // 0x3178
	13'h18bd: q2 = 16'h2068; // 0x317a
	13'h18be: q2 = 16'h0010; // 0x317c
	13'h18bf: q2 = 16'h2028; // 0x317e
	13'h18c0: q2 = 16'h0012; // 0x3180
	13'h18c1: q2 = 16'h90bc; // 0x3182
	13'h18c2: q2 = 16'h0001; // 0x3184
	13'h18c3: q2 = 16'h8072; // 0x3186
	13'h18c4: q2 = 16'he680; // 0x3188
	13'h18c5: q2 = 16'h3680; // 0x318a
	13'h18c6: q2 = 16'h548b; // 0x318c
	13'h18c7: q2 = 16'h206e; // 0x318e
	13'h18c8: q2 = 16'hfff4; // 0x3190
	13'h18c9: q2 = 16'h2068; // 0x3192
	13'h18ca: q2 = 16'h0010; // 0x3194
	13'h18cb: q2 = 16'h2028; // 0x3196
	13'h18cc: q2 = 16'h0012; // 0x3198
	13'h18cd: q2 = 16'h90bc; // 0x319a
	13'h18ce: q2 = 16'h0001; // 0x319c
	13'h18cf: q2 = 16'h8072; // 0x319e
	13'h18d0: q2 = 16'he680; // 0x31a0
	13'h18d1: q2 = 16'he380; // 0x31a2
	13'h18d2: q2 = 16'hd08e; // 0x31a4
	13'h18d3: q2 = 16'h2040; // 0x31a6
	13'h18d4: q2 = 16'h317c; // 0x31a8
	13'h18d5: q2 = 16'h0001; // 0x31aa
	13'h18d6: q2 = 16'hff90; // 0x31ac
	13'h18d7: q2 = 16'h6000; // 0x31ae
	13'h18d8: q2 = 16'hfe3a; // 0x31b0
	13'h18d9: q2 = 16'h7c14; // 0x31b2
	13'h18da: q2 = 16'h41ee; // 0x31b4
	13'h18db: q2 = 16'hffb8; // 0x31b6
	13'h18dc: q2 = 16'h2d48; // 0x31b8
	13'h18dd: q2 = 16'hff8c; // 0x31ba
	13'h18de: q2 = 16'hbc7c; // 0x31bc
	13'h18df: q2 = 16'h002d; // 0x31be
	13'h18e0: q2 = 16'h6e24; // 0x31c0
	13'h18e1: q2 = 16'h206e; // 0x31c2
	13'h18e2: q2 = 16'hff8c; // 0x31c4
	13'h18e3: q2 = 16'h4a50; // 0x31c6
	13'h18e4: q2 = 16'h6614; // 0x31c8
	13'h18e5: q2 = 16'h3686; // 0x31ca
	13'h18e6: q2 = 16'h548b; // 0x31cc
	13'h18e7: q2 = 16'h3006; // 0x31ce
	13'h18e8: q2 = 16'he340; // 0x31d0
	13'h18e9: q2 = 16'h48c0; // 0x31d2
	13'h18ea: q2 = 16'hd08e; // 0x31d4
	13'h18eb: q2 = 16'h2040; // 0x31d6
	13'h18ec: q2 = 16'h317c; // 0x31d8
	13'h18ed: q2 = 16'h0001; // 0x31da
	13'h18ee: q2 = 16'hff90; // 0x31dc
	13'h18ef: q2 = 16'h5246; // 0x31de
	13'h18f0: q2 = 16'h54ae; // 0x31e0
	13'h18f1: q2 = 16'hff8c; // 0x31e2
	13'h18f2: q2 = 16'h60d6; // 0x31e4
	13'h18f3: q2 = 16'h2a7c; // 0x31e6
	13'h18f4: q2 = 16'h0001; // 0x31e8
	13'h18f5: q2 = 16'h86dc; // 0x31ea
	13'h18f6: q2 = 16'h200e; // 0x31ec
	13'h18f7: q2 = 16'hd0bc; // 0x31ee
	13'h18f8: q2 = 16'hffff; // 0x31f0
	13'h18f9: q2 = 16'hff2c; // 0x31f2
	13'h18fa: q2 = 16'h2f00; // 0x31f4
	13'h18fb: q2 = 16'h200b; // 0x31f6
	13'h18fc: q2 = 16'h221f; // 0x31f8
	13'h18fd: q2 = 16'h9081; // 0x31fa
	13'h18fe: q2 = 16'he280; // 0x31fc
	13'h18ff: q2 = 16'h3a00; // 0x31fe
	13'h1900: q2 = 16'h3e39; // 0x3200
	13'h1901: q2 = 16'h0001; // 0x3202
	13'h1902: q2 = 16'h7fa6; // 0x3204
	13'h1903: q2 = 16'h4246; // 0x3206
	13'h1904: q2 = 16'h47ee; // 0x3208
	13'h1905: q2 = 16'hff2c; // 0x320a
	13'h1906: q2 = 16'hbc45; // 0x320c
	13'h1907: q2 = 16'h6c00; // 0x320e
	13'h1908: q2 = 16'h0094; // 0x3210
	13'h1909: q2 = 16'h3013; // 0x3212
	13'h190a: q2 = 16'he340; // 0x3214
	13'h190b: q2 = 16'h48c0; // 0x3216
	13'h190c: q2 = 16'hd08e; // 0x3218
	13'h190d: q2 = 16'h2040; // 0x321a
	13'h190e: q2 = 16'h4a68; // 0x321c
	13'h190f: q2 = 16'hff90; // 0x321e
	13'h1910: q2 = 16'h6700; // 0x3220
	13'h1911: q2 = 16'h007a; // 0x3222
	13'h1912: q2 = 16'h3013; // 0x3224
	13'h1913: q2 = 16'he740; // 0x3226
	13'h1914: q2 = 16'h48c0; // 0x3228
	13'h1915: q2 = 16'h2840; // 0x322a
	13'h1916: q2 = 16'hd9fc; // 0x322c
	13'h1917: q2 = 16'h0001; // 0x322e
	13'h1918: q2 = 16'h8072; // 0x3230
	13'h1919: q2 = 16'h3014; // 0x3232
	13'h191a: q2 = 16'hee40; // 0x3234
	13'h191b: q2 = 16'h5340; // 0x3236
	13'h191c: q2 = 16'h1b40; // 0x3238
	13'h191d: q2 = 16'h0002; // 0x323a
	13'h191e: q2 = 16'h4a47; // 0x323c
	13'h191f: q2 = 16'h6710; // 0x323e
	13'h1920: q2 = 16'h303c; // 0x3240
	13'h1921: q2 = 16'h00ee; // 0x3242
	13'h1922: q2 = 16'h122d; // 0x3244
	13'h1923: q2 = 16'h0002; // 0x3246
	13'h1924: q2 = 16'h4881; // 0x3248
	13'h1925: q2 = 16'h9041; // 0x324a
	13'h1926: q2 = 16'h1b40; // 0x324c
	13'h1927: q2 = 16'h0002; // 0x324e
	13'h1928: q2 = 16'h302c; // 0x3250
	13'h1929: q2 = 16'h0002; // 0x3252
	13'h192a: q2 = 16'hee40; // 0x3254
	13'h192b: q2 = 16'h1b40; // 0x3256
	13'h192c: q2 = 16'h0003; // 0x3258
	13'h192d: q2 = 16'h4a47; // 0x325a
	13'h192e: q2 = 16'h6716; // 0x325c
	13'h192f: q2 = 16'h4a2d; // 0x325e
	13'h1930: q2 = 16'h0003; // 0x3260
	13'h1931: q2 = 16'h6710; // 0x3262
	13'h1932: q2 = 16'h303c; // 0x3264
	13'h1933: q2 = 16'h0112; // 0x3266
	13'h1934: q2 = 16'h122d; // 0x3268
	13'h1935: q2 = 16'h0003; // 0x326a
	13'h1936: q2 = 16'h4881; // 0x326c
	13'h1937: q2 = 16'h9041; // 0x326e
	13'h1938: q2 = 16'h1b40; // 0x3270
	13'h1939: q2 = 16'h0003; // 0x3272
	13'h193a: q2 = 16'h302c; // 0x3274
	13'h193b: q2 = 16'h0006; // 0x3276
	13'h193c: q2 = 16'hc07c; // 0x3278
	13'h193d: q2 = 16'h00ff; // 0x327a
	13'h193e: q2 = 16'h1a80; // 0x327c
	13'h193f: q2 = 16'h4a47; // 0x327e
	13'h1940: q2 = 16'h670c; // 0x3280
	13'h1941: q2 = 16'h1015; // 0x3282
	13'h1942: q2 = 16'h4880; // 0x3284
	13'h1943: q2 = 16'h323c; // 0x3286
	13'h1944: q2 = 16'h00c0; // 0x3288
	13'h1945: q2 = 16'hb340; // 0x328a
	13'h1946: q2 = 16'h1a80; // 0x328c
	13'h1947: q2 = 16'h302c; // 0x328e
	13'h1948: q2 = 16'h0004; // 0x3290
	13'h1949: q2 = 16'hc07c; // 0x3292
	13'h194a: q2 = 16'h00ff; // 0x3294
	13'h194b: q2 = 16'h1b40; // 0x3296
	13'h194c: q2 = 16'h0001; // 0x3298
	13'h194d: q2 = 16'h588d; // 0x329a
	13'h194e: q2 = 16'h5246; // 0x329c
	13'h194f: q2 = 16'h548b; // 0x329e
	13'h1950: q2 = 16'h6000; // 0x32a0
	13'h1951: q2 = 16'hff6a; // 0x32a2
	13'h1952: q2 = 16'h4a9f; // 0x32a4
	13'h1953: q2 = 16'h4cdf; // 0x32a6
	13'h1954: q2 = 16'h38f0; // 0x32a8
	13'h1955: q2 = 16'h4e5e; // 0x32aa
	13'h1956: q2 = 16'h4e75; // 0x32ac
	13'h1957: q2 = 16'h4e56; // 0x32ae
	13'h1958: q2 = 16'h0000; // 0x32b0
	13'h1959: q2 = 16'h48e7; // 0x32b2
	13'h195a: q2 = 16'h0700; // 0x32b4
	13'h195b: q2 = 16'h4247; // 0x32b6
	13'h195c: q2 = 16'hbe7c; // 0x32b8
	13'h195d: q2 = 16'h000a; // 0x32ba
	13'h195e: q2 = 16'h6c00; // 0x32bc
	13'h195f: q2 = 16'h009e; // 0x32be
	13'h1960: q2 = 16'h3007; // 0x32c0
	13'h1961: q2 = 16'he340; // 0x32c2
	13'h1962: q2 = 16'h48c0; // 0x32c4
	13'h1963: q2 = 16'hd0bc; // 0x32c6
	13'h1964: q2 = 16'h0001; // 0x32c8
	13'h1965: q2 = 16'h86b8; // 0x32ca
	13'h1966: q2 = 16'h2040; // 0x32cc
	13'h1967: q2 = 16'h3c10; // 0x32ce
	13'h1968: q2 = 16'h3007; // 0x32d0
	13'h1969: q2 = 16'h6000; // 0x32d2
	13'h196a: q2 = 16'h006e; // 0x32d4
	13'h196b: q2 = 16'h3006; // 0x32d6
	13'h196c: q2 = 16'h5440; // 0x32d8
	13'h196d: q2 = 16'h33c0; // 0x32da
	13'h196e: q2 = 16'h0001; // 0x32dc
	13'h196f: q2 = 16'h757a; // 0x32de
	13'h1970: q2 = 16'h6000; // 0x32e0
	13'h1971: q2 = 16'h0074; // 0x32e2
	13'h1972: q2 = 16'h3006; // 0x32e4
	13'h1973: q2 = 16'h5240; // 0x32e6
	13'h1974: q2 = 16'h33c0; // 0x32e8
	13'h1975: q2 = 16'h0001; // 0x32ea
	13'h1976: q2 = 16'h757e; // 0x32ec
	13'h1977: q2 = 16'h6066; // 0x32ee
	13'h1978: q2 = 16'h3006; // 0x32f0
	13'h1979: q2 = 16'hc1fc; // 0x32f2
	13'h197a: q2 = 16'h0032; // 0x32f4
	13'h197b: q2 = 16'h33c0; // 0x32f6
	13'h197c: q2 = 16'h0001; // 0x32f8
	13'h197d: q2 = 16'h7580; // 0x32fa
	13'h197e: q2 = 16'h6058; // 0x32fc
	13'h197f: q2 = 16'h3006; // 0x32fe
	13'h1980: q2 = 16'hc1fc; // 0x3300
	13'h1981: q2 = 16'h0032; // 0x3302
	13'h1982: q2 = 16'h33c0; // 0x3304
	13'h1983: q2 = 16'h0001; // 0x3306
	13'h1984: q2 = 16'h7582; // 0x3308
	13'h1985: q2 = 16'h604a; // 0x330a
	13'h1986: q2 = 16'h33c6; // 0x330c
	13'h1987: q2 = 16'h0001; // 0x330e
	13'h1988: q2 = 16'h7586; // 0x3310
	13'h1989: q2 = 16'h6042; // 0x3312
	13'h198a: q2 = 16'h33c6; // 0x3314
	13'h198b: q2 = 16'h0001; // 0x3316
	13'h198c: q2 = 16'h7588; // 0x3318
	13'h198d: q2 = 16'h603a; // 0x331a
	13'h198e: q2 = 16'h33c6; // 0x331c
	13'h198f: q2 = 16'h0001; // 0x331e
	13'h1990: q2 = 16'h758a; // 0x3320
	13'h1991: q2 = 16'h6032; // 0x3322
	13'h1992: q2 = 16'h33c6; // 0x3324
	13'h1993: q2 = 16'h0001; // 0x3326
	13'h1994: q2 = 16'h758c; // 0x3328
	13'h1995: q2 = 16'h602a; // 0x332a
	13'h1996: q2 = 16'h33c6; // 0x332c
	13'h1997: q2 = 16'h0001; // 0x332e
	13'h1998: q2 = 16'h758e; // 0x3330
	13'h1999: q2 = 16'h6022; // 0x3332
	13'h199a: q2 = 16'h3006; // 0x3334
	13'h199b: q2 = 16'h5240; // 0x3336
	13'h199c: q2 = 16'h33c0; // 0x3338
	13'h199d: q2 = 16'h0001; // 0x333a
	13'h199e: q2 = 16'h7592; // 0x333c
	13'h199f: q2 = 16'h6016; // 0x333e
	13'h19a0: q2 = 16'h6014; // 0x3340
	13'h19a1: q2 = 16'hb07c; // 0x3342
	13'h19a2: q2 = 16'h0009; // 0x3344
	13'h19a3: q2 = 16'h620e; // 0x3346
	13'h19a4: q2 = 16'he540; // 0x3348
	13'h19a5: q2 = 16'h3040; // 0x334a
	13'h19a6: q2 = 16'hd1fc; // 0x334c
	13'h19a7: q2 = 16'h0000; // 0x334e
	13'h19a8: q2 = 16'hfd26; // 0x3350
	13'h19a9: q2 = 16'h2050; // 0x3352
	13'h19aa: q2 = 16'h4ed0; // 0x3354
	13'h19ab: q2 = 16'h5247; // 0x3356
	13'h19ac: q2 = 16'h6000; // 0x3358
	13'h19ad: q2 = 16'hff5e; // 0x335a
	13'h19ae: q2 = 16'h4a9f; // 0x335c
	13'h19af: q2 = 16'h4cdf; // 0x335e
	13'h19b0: q2 = 16'h00c0; // 0x3360
	13'h19b1: q2 = 16'h4e5e; // 0x3362
	13'h19b2: q2 = 16'h4e75; // 0x3364
	13'h19b3: q2 = 16'h48e7; // 0x3366
	13'h19b4: q2 = 16'h0018; // 0x3368
	13'h19b5: q2 = 16'h701c; // 0x336a
	13'h19b6: q2 = 16'h207c; // 0x336c
	13'h19b7: q2 = 16'h0001; // 0x336e
	13'h19b8: q2 = 16'h7808; // 0x3370
	13'h19b9: q2 = 16'h227c; // 0x3372
	13'h19ba: q2 = 16'h0001; // 0x3374
	13'h19bb: q2 = 16'h7a00; // 0x3376
	13'h19bc: q2 = 16'h247c; // 0x3378
	13'h19bd: q2 = 16'h0001; // 0x337a
	13'h19be: q2 = 16'h77ea; // 0x337c
	13'h19bf: q2 = 16'h267c; // 0x337e
	13'h19c0: q2 = 16'h0000; // 0x3380
	13'h19c1: q2 = 16'hca60; // 0x3382
	13'h19c2: q2 = 16'h287c; // 0x3384
	13'h19c3: q2 = 16'h0000; // 0x3386
	13'h19c4: q2 = 16'hca7e; // 0x3388
	13'h19c5: q2 = 16'h3233; // 0x338a
	13'h19c6: q2 = 16'h0000; // 0x338c
	13'h19c7: q2 = 16'h6d0c; // 0x338e
	13'h19c8: q2 = 16'h42b0; // 0x3390
	13'h19c9: q2 = 16'h1000; // 0x3392
	13'h19ca: q2 = 16'h42b0; // 0x3394
	13'h19cb: q2 = 16'h100c; // 0x3396
	13'h19cc: q2 = 16'h42b0; // 0x3398
	13'h19cd: q2 = 16'h1018; // 0x339a
	13'h19ce: q2 = 16'h3234; // 0x339c
	13'h19cf: q2 = 16'h0000; // 0x339e
	13'h19d0: q2 = 16'h42b0; // 0x33a0
	13'h19d1: q2 = 16'h1000; // 0x33a2
	13'h19d2: q2 = 16'h4271; // 0x33a4
	13'h19d3: q2 = 16'h0000; // 0x33a6
	13'h19d4: q2 = 16'h4272; // 0x33a8
	13'h19d5: q2 = 16'h0000; // 0x33aa
	13'h19d6: q2 = 16'h5540; // 0x33ac
	13'h19d7: q2 = 16'h6cda; // 0x33ae
	13'h19d8: q2 = 16'h33fc; // 0x33b0
	13'h19d9: q2 = 16'h0001; // 0x33b2
	13'h19da: q2 = 16'h0001; // 0x33b4
	13'h19db: q2 = 16'h7a3c; // 0x33b6
	13'h19dc: q2 = 16'h33fc; // 0x33b8
	13'h19dd: q2 = 16'hffff; // 0x33ba
	13'h19de: q2 = 16'h0001; // 0x33bc
	13'h19df: q2 = 16'h7b9c; // 0x33be
	13'h19e0: q2 = 16'h4cdf; // 0x33c0
	13'h19e1: q2 = 16'h1800; // 0x33c2
	13'h19e2: q2 = 16'h4e75; // 0x33c4
	13'h19e3: q2 = 16'h4e56; // 0x33c6
	13'h19e4: q2 = 16'hfff8; // 0x33c8
	13'h19e5: q2 = 16'h48e7; // 0x33ca
	13'h19e6: q2 = 16'h0704; // 0x33cc
	13'h19e7: q2 = 16'h2a79; // 0x33ce
	13'h19e8: q2 = 16'h0001; // 0x33d0
	13'h19e9: q2 = 16'h7fb8; // 0x33d2
	13'h19ea: q2 = 16'h3ebc; // 0x33d4
	13'h19eb: q2 = 16'h001b; // 0x33d6
	13'h19ec: q2 = 16'h4eb9; // 0x33d8
	13'h19ed: q2 = 16'h0000; // 0x33da
	13'h19ee: q2 = 16'h8a22; // 0x33dc
	13'h19ef: q2 = 16'h4a79; // 0x33de
	13'h19f0: q2 = 16'h0001; // 0x33e0
	13'h19f1: q2 = 16'h7fc6; // 0x33e2
	13'h19f2: q2 = 16'h6720; // 0x33e4
	13'h19f3: q2 = 16'h3ebc; // 0x33e6
	13'h19f4: q2 = 16'h0029; // 0x33e8
	13'h19f5: q2 = 16'h4267; // 0x33ea
	13'h19f6: q2 = 16'h3f3c; // 0x33ec
	13'h19f7: q2 = 16'hffe1; // 0x33ee
	13'h19f8: q2 = 16'h3f3c; // 0x33f0
	13'h19f9: q2 = 16'h0004; // 0x33f2
	13'h19fa: q2 = 16'h2f3c; // 0x33f4
	13'h19fb: q2 = 16'h0000; // 0x33f6
	13'h19fc: q2 = 16'hb488; // 0x33f8
	13'h19fd: q2 = 16'h4eb9; // 0x33fa
	13'h19fe: q2 = 16'h0000; // 0x33fc
	13'h19ff: q2 = 16'h026c; // 0x33fe
	13'h1a00: q2 = 16'hdefc; // 0x3400
	13'h1a01: q2 = 16'h000a; // 0x3402
	13'h1a02: q2 = 16'h600a; // 0x3404
	13'h1a03: q2 = 16'h3ebc; // 0x3406
	13'h1a04: q2 = 16'h000b; // 0x3408
	13'h1a05: q2 = 16'h4eb9; // 0x340a
	13'h1a06: q2 = 16'h0000; // 0x340c
	13'h1a07: q2 = 16'h549c; // 0x340e
	13'h1a08: q2 = 16'h4eb9; // 0x3410
	13'h1a09: q2 = 16'h0000; // 0x3412
	13'h1a0a: q2 = 16'h8a92; // 0x3414
	13'h1a0b: q2 = 16'h200e; // 0x3416
	13'h1a0c: q2 = 16'hd0bc; // 0x3418
	13'h1a0d: q2 = 16'hffff; // 0x341a
	13'h1a0e: q2 = 16'hfff8; // 0x341c
	13'h1a0f: q2 = 16'h2e80; // 0x341e
	13'h1a10: q2 = 16'h3f15; // 0x3420
	13'h1a11: q2 = 16'h4eb9; // 0x3422
	13'h1a12: q2 = 16'h0000; // 0x3424
	13'h1a13: q2 = 16'h0828; // 0x3426
	13'h1a14: q2 = 16'h4a5f; // 0x3428
	13'h1a15: q2 = 16'h0c79; // 0x342a
	13'h1a16: q2 = 16'h0003; // 0x342c
	13'h1a17: q2 = 16'h0001; // 0x342e
	13'h1a18: q2 = 16'h758c; // 0x3430
	13'h1a19: q2 = 16'h6604; // 0x3432
	13'h1a1a: q2 = 16'h7c07; // 0x3434
	13'h1a1b: q2 = 16'h6002; // 0x3436
	13'h1a1c: q2 = 16'h7c06; // 0x3438
	13'h1a1d: q2 = 16'h4247; // 0x343a
	13'h1a1e: q2 = 16'h200e; // 0x343c
	13'h1a1f: q2 = 16'hd0bc; // 0x343e
	13'h1a20: q2 = 16'hffff; // 0x3440
	13'h1a21: q2 = 16'hfff8; // 0x3442
	13'h1a22: q2 = 16'h2e80; // 0x3444
	13'h1a23: q2 = 16'h4eb9; // 0x3446
	13'h1a24: q2 = 16'h0000; // 0x3448
	13'h1a25: q2 = 16'h072e; // 0x344a
	13'h1a26: q2 = 16'hb047; // 0x344c
	13'h1a27: q2 = 16'h6f2e; // 0x344e
	13'h1a28: q2 = 16'h3e87; // 0x3450
	13'h1a29: q2 = 16'h0657; // 0x3452
	13'h1a2a: q2 = 16'h0022; // 0x3454
	13'h1a2b: q2 = 16'h3207; // 0x3456
	13'h1a2c: q2 = 16'h48c1; // 0x3458
	13'h1a2d: q2 = 16'h200e; // 0x345a
	13'h1a2e: q2 = 16'hd081; // 0x345c
	13'h1a2f: q2 = 16'h2040; // 0x345e
	13'h1a30: q2 = 16'h1028; // 0x3460
	13'h1a31: q2 = 16'hfff8; // 0x3462
	13'h1a32: q2 = 16'h4880; // 0x3464
	13'h1a33: q2 = 16'h3f00; // 0x3466
	13'h1a34: q2 = 16'h3f3c; // 0x3468
	13'h1a35: q2 = 16'h0004; // 0x346a
	13'h1a36: q2 = 16'h3f07; // 0x346c
	13'h1a37: q2 = 16'h3006; // 0x346e
	13'h1a38: q2 = 16'hd157; // 0x3470
	13'h1a39: q2 = 16'h4eb9; // 0x3472
	13'h1a3a: q2 = 16'h0000; // 0x3474
	13'h1a3b: q2 = 16'h3d18; // 0x3476
	13'h1a3c: q2 = 16'h5c4f; // 0x3478
	13'h1a3d: q2 = 16'h5247; // 0x347a
	13'h1a3e: q2 = 16'h60be; // 0x347c
	13'h1a3f: q2 = 16'h4a9f; // 0x347e
	13'h1a40: q2 = 16'h4cdf; // 0x3480
	13'h1a41: q2 = 16'h20c0; // 0x3482
	13'h1a42: q2 = 16'h4e5e; // 0x3484
	13'h1a43: q2 = 16'h4e75; // 0x3486
	13'h1a44: q2 = 16'h234d; // 0x3488
	13'h1a45: q2 = 16'h434d; // 0x348a
	13'h1a46: q2 = 16'h4c58; // 0x348c
	13'h1a47: q2 = 16'h5858; // 0x348e
	13'h1a48: q2 = 16'h4949; // 0x3490
	13'h1a49: q2 = 16'h2041; // 0x3492
	13'h1a4a: q2 = 16'h5441; // 0x3494
	13'h1a4b: q2 = 16'h5249; // 0x3496
	13'h1a4c: q2 = 16'h0000; // 0x3498
	13'h1a4d: q2 = 16'h4e56; // 0x349a
	13'h1a4e: q2 = 16'hff94; // 0x349c
	13'h1a4f: q2 = 16'h48e7; // 0x349e
	13'h1a50: q2 = 16'h1f1c; // 0x34a0
	13'h1a51: q2 = 16'h4eb9; // 0x34a2
	13'h1a52: q2 = 16'h0000; // 0x34a4
	13'h1a53: q2 = 16'h0226; // 0x34a6
	13'h1a54: q2 = 16'h4247; // 0x34a8
	13'h1a55: q2 = 16'hbe7c; // 0x34aa
	13'h1a56: q2 = 16'h0020; // 0x34ac
	13'h1a57: q2 = 16'h6c2c; // 0x34ae
	13'h1a58: q2 = 16'h7c1f; // 0x34b0
	13'h1a59: q2 = 16'hbc7c; // 0x34b2
	13'h1a5a: q2 = 16'h0019; // 0x34b4
	13'h1a5b: q2 = 16'h6d20; // 0x34b6
	13'h1a5c: q2 = 16'h3a06; // 0x34b8
	13'h1a5d: q2 = 16'heb45; // 0x34ba
	13'h1a5e: q2 = 16'hda47; // 0x34bc
	13'h1a5f: q2 = 16'hda7c; // 0x34be
	13'h1a60: q2 = 16'hfe00; // 0x34c0
	13'h1a61: q2 = 16'h3ebc; // 0x34c2
	13'h1a62: q2 = 16'h002c; // 0x34c4
	13'h1a63: q2 = 16'h3f05; // 0x34c6
	13'h1a64: q2 = 16'h3f06; // 0x34c8
	13'h1a65: q2 = 16'h3f07; // 0x34ca
	13'h1a66: q2 = 16'h4eb9; // 0x34cc
	13'h1a67: q2 = 16'h0000; // 0x34ce
	13'h1a68: q2 = 16'h3d18; // 0x34d0
	13'h1a69: q2 = 16'h5c4f; // 0x34d2
	13'h1a6a: q2 = 16'h5346; // 0x34d4
	13'h1a6b: q2 = 16'h60da; // 0x34d6
	13'h1a6c: q2 = 16'h5247; // 0x34d8
	13'h1a6d: q2 = 16'h60ce; // 0x34da
	13'h1a6e: q2 = 16'h3ebc; // 0x34dc
	13'h1a6f: q2 = 16'h003e; // 0x34de
	13'h1a70: q2 = 16'h4267; // 0x34e0
	13'h1a71: q2 = 16'h3f3c; // 0x34e2
	13'h1a72: q2 = 16'h0064; // 0x34e4
	13'h1a73: q2 = 16'h3f3c; // 0x34e6
	13'h1a74: q2 = 16'h0017; // 0x34e8
	13'h1a75: q2 = 16'h2f3c; // 0x34ea
	13'h1a76: q2 = 16'h0000; // 0x34ec
	13'h1a77: q2 = 16'hfe26; // 0x34ee
	13'h1a78: q2 = 16'h4eb9; // 0x34f0
	13'h1a79: q2 = 16'h0000; // 0x34f2
	13'h1a7a: q2 = 16'h026c; // 0x34f4
	13'h1a7b: q2 = 16'hdefc; // 0x34f6
	13'h1a7c: q2 = 16'h000a; // 0x34f8
	13'h1a7d: q2 = 16'h267c; // 0x34fa
	13'h1a7e: q2 = 16'h0001; // 0x34fc
	13'h1a7f: q2 = 16'h75e8; // 0x34fe
	13'h1a80: q2 = 16'h2d7c; // 0x3500
	13'h1a81: q2 = 16'h0001; // 0x3502
	13'h1a82: q2 = 16'h7ba8; // 0x3504
	13'h1a83: q2 = 16'hffdc; // 0x3506
	13'h1a84: q2 = 16'h2a7c; // 0x3508
	13'h1a85: q2 = 16'h0000; // 0x350a
	13'h1a86: q2 = 16'hfe06; // 0x350c
	13'h1a87: q2 = 16'h287c; // 0x350e
	13'h1a88: q2 = 16'h0000; // 0x3510
	13'h1a89: q2 = 16'hfe16; // 0x3512
	13'h1a8a: q2 = 16'h4247; // 0x3514
	13'h1a8b: q2 = 16'hbe7c; // 0x3516
	13'h1a8c: q2 = 16'h000f; // 0x3518
	13'h1a8d: q2 = 16'h6c00; // 0x351a
	13'h1a8e: q2 = 16'h023e; // 0x351c
	13'h1a8f: q2 = 16'h4246; // 0x351e
	13'h1a90: q2 = 16'hbc7c; // 0x3520
	13'h1a91: q2 = 16'h0003; // 0x3522
	13'h1a92: q2 = 16'h6c32; // 0x3524
	13'h1a93: q2 = 16'h202e; // 0x3526
	13'h1a94: q2 = 16'hffdc; // 0x3528
	13'h1a95: q2 = 16'h2040; // 0x352a
	13'h1a96: q2 = 16'h1a10; // 0x352c
	13'h1a97: q2 = 16'h4885; // 0x352e
	13'h1a98: q2 = 16'h3e87; // 0x3530
	13'h1a99: q2 = 16'h0657; // 0x3532
	13'h1a9a: q2 = 16'h002d; // 0x3534
	13'h1a9b: q2 = 16'h3f05; // 0x3536
	13'h1a9c: q2 = 16'h1014; // 0x3538
	13'h1a9d: q2 = 16'h4880; // 0x353a
	13'h1a9e: q2 = 16'h3f00; // 0x353c
	13'h1a9f: q2 = 16'h1015; // 0x353e
	13'h1aa0: q2 = 16'h4880; // 0x3540
	13'h1aa1: q2 = 16'h3f00; // 0x3542
	13'h1aa2: q2 = 16'h3006; // 0x3544
	13'h1aa3: q2 = 16'hd157; // 0x3546
	13'h1aa4: q2 = 16'h4eb9; // 0x3548
	13'h1aa5: q2 = 16'h0000; // 0x354a
	13'h1aa6: q2 = 16'h3d18; // 0x354c
	13'h1aa7: q2 = 16'h5c4f; // 0x354e
	13'h1aa8: q2 = 16'h5246; // 0x3550
	13'h1aa9: q2 = 16'h52ae; // 0x3552
	13'h1aaa: q2 = 16'hffdc; // 0x3554
	13'h1aab: q2 = 16'h60c8; // 0x3556
	13'h1aac: q2 = 16'h422e; // 0x3558
	13'h1aad: q2 = 16'hfff4; // 0x355a
	13'h1aae: q2 = 16'h200e; // 0x355c
	13'h1aaf: q2 = 16'hd0bc; // 0x355e
	13'h1ab0: q2 = 16'hffff; // 0x3560
	13'h1ab1: q2 = 16'hffe8; // 0x3562
	13'h1ab2: q2 = 16'h2e80; // 0x3564
	13'h1ab3: q2 = 16'h3007; // 0x3566
	13'h1ab4: q2 = 16'he540; // 0x3568
	13'h1ab5: q2 = 16'h48c0; // 0x356a
	13'h1ab6: q2 = 16'hd0bc; // 0x356c
	13'h1ab7: q2 = 16'h0001; // 0x356e
	13'h1ab8: q2 = 16'h7f64; // 0x3570
	13'h1ab9: q2 = 16'h2040; // 0x3572
	13'h1aba: q2 = 16'h2f10; // 0x3574
	13'h1abb: q2 = 16'h4eb9; // 0x3576
	13'h1abc: q2 = 16'h0000; // 0x3578
	13'h1abd: q2 = 16'h0892; // 0x357a
	13'h1abe: q2 = 16'h4a9f; // 0x357c
	13'h1abf: q2 = 16'hbe7c; // 0x357e
	13'h1ac0: q2 = 16'h0003; // 0x3580
	13'h1ac1: q2 = 16'h6c18; // 0x3582
	13'h1ac2: q2 = 16'h2ebc; // 0x3584
	13'h1ac3: q2 = 16'h0000; // 0x3586
	13'h1ac4: q2 = 16'hfe3d; // 0x3588
	13'h1ac5: q2 = 16'h200e; // 0x358a
	13'h1ac6: q2 = 16'hd0bc; // 0x358c
	13'h1ac7: q2 = 16'hffff; // 0x358e
	13'h1ac8: q2 = 16'hfff4; // 0x3590
	13'h1ac9: q2 = 16'h2f00; // 0x3592
	13'h1aca: q2 = 16'h4eb9; // 0x3594
	13'h1acb: q2 = 16'h0000; // 0x3596
	13'h1acc: q2 = 16'h0770; // 0x3598
	13'h1acd: q2 = 16'h4a9f; // 0x359a
	13'h1ace: q2 = 16'h200e; // 0x359c
	13'h1acf: q2 = 16'hd0bc; // 0x359e
	13'h1ad0: q2 = 16'hffff; // 0x35a0
	13'h1ad1: q2 = 16'hffe8; // 0x35a2
	13'h1ad2: q2 = 16'h2e80; // 0x35a4
	13'h1ad3: q2 = 16'h4eb9; // 0x35a6
	13'h1ad4: q2 = 16'h0000; // 0x35a8
	13'h1ad5: q2 = 16'h072e; // 0x35aa
	13'h1ad6: q2 = 16'h3c00; // 0x35ac
	13'h1ad7: q2 = 16'hbc7c; // 0x35ae
	13'h1ad8: q2 = 16'h0008; // 0x35b0
	13'h1ad9: q2 = 16'h6c1c; // 0x35b2
	13'h1ada: q2 = 16'h2ebc; // 0x35b4
	13'h1adb: q2 = 16'h0000; // 0x35b6
	13'h1adc: q2 = 16'hfe3f; // 0x35b8
	13'h1add: q2 = 16'h200e; // 0x35ba
	13'h1ade: q2 = 16'hd0bc; // 0x35bc
	13'h1adf: q2 = 16'hffff; // 0x35be
	13'h1ae0: q2 = 16'hfff4; // 0x35c0
	13'h1ae1: q2 = 16'h2f00; // 0x35c2
	13'h1ae2: q2 = 16'h4eb9; // 0x35c4
	13'h1ae3: q2 = 16'h0000; // 0x35c6
	13'h1ae4: q2 = 16'h0770; // 0x35c8
	13'h1ae5: q2 = 16'h4a9f; // 0x35ca
	13'h1ae6: q2 = 16'h5246; // 0x35cc
	13'h1ae7: q2 = 16'h60de; // 0x35ce
	13'h1ae8: q2 = 16'h200e; // 0x35d0
	13'h1ae9: q2 = 16'hd0bc; // 0x35d2
	13'h1aea: q2 = 16'hffff; // 0x35d4
	13'h1aeb: q2 = 16'hffe8; // 0x35d6
	13'h1aec: q2 = 16'h2e80; // 0x35d8
	13'h1aed: q2 = 16'h200e; // 0x35da
	13'h1aee: q2 = 16'hd0bc; // 0x35dc
	13'h1aef: q2 = 16'hffff; // 0x35de
	13'h1af0: q2 = 16'hfff4; // 0x35e0
	13'h1af1: q2 = 16'h2f00; // 0x35e2
	13'h1af2: q2 = 16'h4eb9; // 0x35e4
	13'h1af3: q2 = 16'h0000; // 0x35e6
	13'h1af4: q2 = 16'h0770; // 0x35e8
	13'h1af5: q2 = 16'h4a9f; // 0x35ea
	13'h1af6: q2 = 16'h2ebc; // 0x35ec
	13'h1af7: q2 = 16'h0000; // 0x35ee
	13'h1af8: q2 = 16'hfe41; // 0x35f0
	13'h1af9: q2 = 16'h200e; // 0x35f2
	13'h1afa: q2 = 16'hd0bc; // 0x35f4
	13'h1afb: q2 = 16'hffff; // 0x35f6
	13'h1afc: q2 = 16'hfff4; // 0x35f8
	13'h1afd: q2 = 16'h2f00; // 0x35fa
	13'h1afe: q2 = 16'h4eb9; // 0x35fc
	13'h1aff: q2 = 16'h0000; // 0x35fe
	13'h1b00: q2 = 16'h0770; // 0x3600
	13'h1b01: q2 = 16'h4a9f; // 0x3602
	13'h1b02: q2 = 16'h4246; // 0x3604
	13'h1b03: q2 = 16'h200e; // 0x3606
	13'h1b04: q2 = 16'hd0bc; // 0x3608
	13'h1b05: q2 = 16'hffff; // 0x360a
	13'h1b06: q2 = 16'hfff4; // 0x360c
	13'h1b07: q2 = 16'h2e80; // 0x360e
	13'h1b08: q2 = 16'h4eb9; // 0x3610
	13'h1b09: q2 = 16'h0000; // 0x3612
	13'h1b0a: q2 = 16'h072e; // 0x3614
	13'h1b0b: q2 = 16'hb046; // 0x3616
	13'h1b0c: q2 = 16'h6f36; // 0x3618
	13'h1b0d: q2 = 16'h3e87; // 0x361a
	13'h1b0e: q2 = 16'h0657; // 0x361c
	13'h1b0f: q2 = 16'h002d; // 0x361e
	13'h1b10: q2 = 16'h3206; // 0x3620
	13'h1b11: q2 = 16'h48c1; // 0x3622
	13'h1b12: q2 = 16'h200e; // 0x3624
	13'h1b13: q2 = 16'hd081; // 0x3626
	13'h1b14: q2 = 16'h2040; // 0x3628
	13'h1b15: q2 = 16'h1028; // 0x362a
	13'h1b16: q2 = 16'hfff4; // 0x362c
	13'h1b17: q2 = 16'h4880; // 0x362e
	13'h1b18: q2 = 16'h3f00; // 0x3630
	13'h1b19: q2 = 16'h1014; // 0x3632
	13'h1b1a: q2 = 16'h4880; // 0x3634
	13'h1b1b: q2 = 16'h3f00; // 0x3636
	13'h1b1c: q2 = 16'h1015; // 0x3638
	13'h1b1d: q2 = 16'h4880; // 0x363a
	13'h1b1e: q2 = 16'h3f00; // 0x363c
	13'h1b1f: q2 = 16'h3006; // 0x363e
	13'h1b20: q2 = 16'hd157; // 0x3640
	13'h1b21: q2 = 16'h5657; // 0x3642
	13'h1b22: q2 = 16'h4eb9; // 0x3644
	13'h1b23: q2 = 16'h0000; // 0x3646
	13'h1b24: q2 = 16'h3d18; // 0x3648
	13'h1b25: q2 = 16'h5c4f; // 0x364a
	13'h1b26: q2 = 16'h5246; // 0x364c
	13'h1b27: q2 = 16'h60b6; // 0x364e
	13'h1b28: q2 = 16'h3e87; // 0x3650
	13'h1b29: q2 = 16'h5257; // 0x3652
	13'h1b2a: q2 = 16'h200e; // 0x3654
	13'h1b2b: q2 = 16'hd0bc; // 0x3656
	13'h1b2c: q2 = 16'hffff; // 0x3658
	13'h1b2d: q2 = 16'hffe2; // 0x365a
	13'h1b2e: q2 = 16'h2f00; // 0x365c
	13'h1b2f: q2 = 16'h200e; // 0x365e
	13'h1b30: q2 = 16'hd0bc; // 0x3660
	13'h1b31: q2 = 16'hffff; // 0x3662
	13'h1b32: q2 = 16'hffe0; // 0x3664
	13'h1b33: q2 = 16'h2f00; // 0x3666
	13'h1b34: q2 = 16'h3007; // 0x3668
	13'h1b35: q2 = 16'he340; // 0x366a
	13'h1b36: q2 = 16'h48c0; // 0x366c
	13'h1b37: q2 = 16'hd0bc; // 0x366e
	13'h1b38: q2 = 16'h0001; // 0x3670
	13'h1b39: q2 = 16'h7efe; // 0x3672
	13'h1b3a: q2 = 16'h2040; // 0x3674
	13'h1b3b: q2 = 16'h3f10; // 0x3676
	13'h1b3c: q2 = 16'h4eb9; // 0x3678
	13'h1b3d: q2 = 16'h0000; // 0x367a
	13'h1b3e: q2 = 16'h1402; // 0x367c
	13'h1b3f: q2 = 16'hdefc; // 0x367e
	13'h1b40: q2 = 16'h000a; // 0x3680
	13'h1b41: q2 = 16'h0c6e; // 0x3682
	13'h1b42: q2 = 16'h0001; // 0x3684
	13'h1b43: q2 = 16'hffe0; // 0x3686
	13'h1b44: q2 = 16'h6606; // 0x3688
	13'h1b45: q2 = 16'h3a3c; // 0x368a
	13'h1b46: q2 = 16'h00e9; // 0x368c
	13'h1b47: q2 = 16'h6012; // 0x368e
	13'h1b48: q2 = 16'h0c6e; // 0x3690
	13'h1b49: q2 = 16'h0002; // 0x3692
	13'h1b4a: q2 = 16'hffe0; // 0x3694
	13'h1b4b: q2 = 16'h6606; // 0x3696
	13'h1b4c: q2 = 16'h3a3c; // 0x3698
	13'h1b4d: q2 = 16'h00e1; // 0x369a
	13'h1b4e: q2 = 16'h6004; // 0x369c
	13'h1b4f: q2 = 16'h3a3c; // 0x369e
	13'h1b50: q2 = 16'h00d9; // 0x36a0
	13'h1b51: q2 = 16'h1c15; // 0x36a2
	13'h1b52: q2 = 16'h4886; // 0x36a4
	13'h1b53: q2 = 16'hdc7c; // 0x36a6
	13'h1b54: q2 = 16'h000e; // 0x36a8
	13'h1b55: q2 = 16'hbe7c; // 0x36aa
	13'h1b56: q2 = 16'h0003; // 0x36ac
	13'h1b57: q2 = 16'h6c02; // 0x36ae
	13'h1b58: q2 = 16'h5246; // 0x36b0
	13'h1b59: q2 = 16'h3e87; // 0x36b2
	13'h1b5a: q2 = 16'h5257; // 0x36b4
	13'h1b5b: q2 = 16'h3f05; // 0x36b6
	13'h1b5c: q2 = 16'h1014; // 0x36b8
	13'h1b5d: q2 = 16'h4880; // 0x36ba
	13'h1b5e: q2 = 16'h3f00; // 0x36bc
	13'h1b5f: q2 = 16'h3f06; // 0x36be
	13'h1b60: q2 = 16'h4eb9; // 0x36c0
	13'h1b61: q2 = 16'h0000; // 0x36c2
	13'h1b62: q2 = 16'h3d18; // 0x36c4
	13'h1b63: q2 = 16'h5c4f; // 0x36c6
	13'h1b64: q2 = 16'h3807; // 0x36c8
	13'h1b65: q2 = 16'hd87c; // 0x36ca
	13'h1b66: q2 = 16'h0010; // 0x36cc
	13'h1b67: q2 = 16'he544; // 0x36ce
	13'h1b68: q2 = 16'h3004; // 0x36d0
	13'h1b69: q2 = 16'he340; // 0x36d2
	13'h1b6a: q2 = 16'h48c0; // 0x36d4
	13'h1b6b: q2 = 16'hd08b; // 0x36d6
	13'h1b6c: q2 = 16'h2040; // 0x36d8
	13'h1b6d: q2 = 16'h316e; // 0x36da
	13'h1b6e: q2 = 16'hffe2; // 0x36dc
	13'h1b6f: q2 = 16'h0002; // 0x36de
	13'h1b70: q2 = 16'h3004; // 0x36e0
	13'h1b71: q2 = 16'he340; // 0x36e2
	13'h1b72: q2 = 16'h48c0; // 0x36e4
	13'h1b73: q2 = 16'hd08b; // 0x36e6
	13'h1b74: q2 = 16'h2040; // 0x36e8
	13'h1b75: q2 = 16'h317c; // 0x36ea
	13'h1b76: q2 = 16'h0013; // 0x36ec
	13'h1b77: q2 = 16'h0004; // 0x36ee
	13'h1b78: q2 = 16'h3004; // 0x36f0
	13'h1b79: q2 = 16'he340; // 0x36f2
	13'h1b7a: q2 = 16'h48c0; // 0x36f4
	13'h1b7b: q2 = 16'hd08b; // 0x36f6
	13'h1b7c: q2 = 16'h2040; // 0x36f8
	13'h1b7d: q2 = 16'h317c; // 0x36fa
	13'h1b7e: q2 = 16'h001d; // 0x36fc
	13'h1b7f: q2 = 16'h0006; // 0x36fe
	13'h1b80: q2 = 16'h3ebc; // 0x3700
	13'h1b81: q2 = 16'h000a; // 0x3702
	13'h1b82: q2 = 16'h4267; // 0x3704
	13'h1b83: q2 = 16'h4eb9; // 0x3706
	13'h1b84: q2 = 16'h0000; // 0x3708
	13'h1b85: q2 = 16'h8e6c; // 0x370a
	13'h1b86: q2 = 16'h4a5f; // 0x370c
	13'h1b87: q2 = 16'h3207; // 0x370e
	13'h1b88: q2 = 16'he341; // 0x3710
	13'h1b89: q2 = 16'h48c1; // 0x3712
	13'h1b8a: q2 = 16'hd28e; // 0x3714
	13'h1b8b: q2 = 16'h2241; // 0x3716
	13'h1b8c: q2 = 16'h3340; // 0x3718
	13'h1b8d: q2 = 16'hff9e; // 0x371a
	13'h1b8e: q2 = 16'h3004; // 0x371c
	13'h1b8f: q2 = 16'he440; // 0x371e
	13'h1b90: q2 = 16'h3e80; // 0x3720
	13'h1b91: q2 = 16'h3007; // 0x3722
	13'h1b92: q2 = 16'he340; // 0x3724
	13'h1b93: q2 = 16'h48c0; // 0x3726
	13'h1b94: q2 = 16'hd08e; // 0x3728
	13'h1b95: q2 = 16'h2040; // 0x372a
	13'h1b96: q2 = 16'h3028; // 0x372c
	13'h1b97: q2 = 16'hff9e; // 0x372e
	13'h1b98: q2 = 16'he340; // 0x3730
	13'h1b99: q2 = 16'h48c0; // 0x3732
	13'h1b9a: q2 = 16'hd0bc; // 0x3734
	13'h1b9b: q2 = 16'h0000; // 0x3736
	13'h1b9c: q2 = 16'hca9c; // 0x3738
	13'h1b9d: q2 = 16'h2040; // 0x373a
	13'h1b9e: q2 = 16'h3f10; // 0x373c
	13'h1b9f: q2 = 16'h1014; // 0x373e
	13'h1ba0: q2 = 16'h4880; // 0x3740
	13'h1ba1: q2 = 16'h3f00; // 0x3742
	13'h1ba2: q2 = 16'h5357; // 0x3744
	13'h1ba3: q2 = 16'h3f06; // 0x3746
	13'h1ba4: q2 = 16'h4eb9; // 0x3748
	13'h1ba5: q2 = 16'h0000; // 0x374a
	13'h1ba6: q2 = 16'h3d18; // 0x374c
	13'h1ba7: q2 = 16'h5c4f; // 0x374e
	13'h1ba8: q2 = 16'h5247; // 0x3750
	13'h1ba9: q2 = 16'h528d; // 0x3752
	13'h1baa: q2 = 16'h528c; // 0x3754
	13'h1bab: q2 = 16'h6000; // 0x3756
	13'h1bac: q2 = 16'hfdbe; // 0x3758
	13'h1bad: q2 = 16'h3d7c; // 0x375a
	13'h1bae: q2 = 16'h0002; // 0x375c
	13'h1baf: q2 = 16'hffda; // 0x375e
	13'h1bb0: q2 = 16'h4247; // 0x3760
	13'h1bb1: q2 = 16'hbe7c; // 0x3762
	13'h1bb2: q2 = 16'h000f; // 0x3764
	13'h1bb3: q2 = 16'h6c1c; // 0x3766
	13'h1bb4: q2 = 16'h3007; // 0x3768
	13'h1bb5: q2 = 16'he340; // 0x376a
	13'h1bb6: q2 = 16'h48c0; // 0x376c
	13'h1bb7: q2 = 16'hd08e; // 0x376e
	13'h1bb8: q2 = 16'h2040; // 0x3770
	13'h1bb9: q2 = 16'h3179; // 0x3772
	13'h1bba: q2 = 16'h0000; // 0x3774
	13'h1bbb: q2 = 16'hcab2; // 0x3776
	13'h1bbc: q2 = 16'hffbc; // 0x3778
	13'h1bbd: q2 = 16'h3d7c; // 0x377a
	13'h1bbe: q2 = 16'h0006; // 0x377c
	13'h1bbf: q2 = 16'hff9c; // 0x377e
	13'h1bc0: q2 = 16'h5247; // 0x3780
	13'h1bc1: q2 = 16'h60de; // 0x3782
	13'h1bc2: q2 = 16'h23fc; // 0x3784
	13'h1bc3: q2 = 16'h0000; // 0x3786
	13'h1bc4: q2 = 16'h0002; // 0x3788
	13'h1bc5: q2 = 16'h0001; // 0x378a
	13'h1bc6: q2 = 16'h7fc2; // 0x378c
	13'h1bc7: q2 = 16'h536e; // 0x378e
	13'h1bc8: q2 = 16'hffda; // 0x3790
	13'h1bc9: q2 = 16'h4a6e; // 0x3792
	13'h1bca: q2 = 16'hffda; // 0x3794
	13'h1bcb: q2 = 16'h6600; // 0x3796
	13'h1bcc: q2 = 16'h00a2; // 0x3798
	13'h1bcd: q2 = 16'h4246; // 0x379a
	13'h1bce: q2 = 16'hbc7c; // 0x379c
	13'h1bcf: q2 = 16'h0004; // 0x379e
	13'h1bd0: q2 = 16'h6c1e; // 0x37a0
	13'h1bd1: q2 = 16'h3006; // 0x37a2
	13'h1bd2: q2 = 16'he340; // 0x37a4
	13'h1bd3: q2 = 16'h48c0; // 0x37a6
	13'h1bd4: q2 = 16'hd08e; // 0x37a8
	13'h1bd5: q2 = 16'h2040; // 0x37aa
	13'h1bd6: q2 = 16'h3206; // 0x37ac
	13'h1bd7: q2 = 16'he341; // 0x37ae
	13'h1bd8: q2 = 16'h48c1; // 0x37b0
	13'h1bd9: q2 = 16'hd28b; // 0x37b2
	13'h1bda: q2 = 16'h2241; // 0x37b4
	13'h1bdb: q2 = 16'h3169; // 0x37b6
	13'h1bdc: q2 = 16'h0168; // 0x37b8
	13'h1bdd: q2 = 16'hff94; // 0x37ba
	13'h1bde: q2 = 16'h5246; // 0x37bc
	13'h1bdf: q2 = 16'h60dc; // 0x37be
	13'h1be0: q2 = 16'h7e2d; // 0x37c0
	13'h1be1: q2 = 16'hbe7c; // 0x37c2
	13'h1be2: q2 = 16'h003f; // 0x37c4
	13'h1be3: q2 = 16'h6c3c; // 0x37c6
	13'h1be4: q2 = 16'h4246; // 0x37c8
	13'h1be5: q2 = 16'hbc7c; // 0x37ca
	13'h1be6: q2 = 16'h0004; // 0x37cc
	13'h1be7: q2 = 16'h6c30; // 0x37ce
	13'h1be8: q2 = 16'h3006; // 0x37d0
	13'h1be9: q2 = 16'he340; // 0x37d2
	13'h1bea: q2 = 16'h48c0; // 0x37d4
	13'h1beb: q2 = 16'h2f00; // 0x37d6
	13'h1bec: q2 = 16'h3007; // 0x37d8
	13'h1bed: q2 = 16'he740; // 0x37da
	13'h1bee: q2 = 16'h48c0; // 0x37dc
	13'h1bef: q2 = 16'h221f; // 0x37de
	13'h1bf0: q2 = 16'hd081; // 0x37e0
	13'h1bf1: q2 = 16'hd08b; // 0x37e2
	13'h1bf2: q2 = 16'h2040; // 0x37e4
	13'h1bf3: q2 = 16'h3206; // 0x37e6
	13'h1bf4: q2 = 16'he341; // 0x37e8
	13'h1bf5: q2 = 16'h48c1; // 0x37ea
	13'h1bf6: q2 = 16'h2241; // 0x37ec
	13'h1bf7: q2 = 16'h3407; // 0x37ee
	13'h1bf8: q2 = 16'he742; // 0x37f0
	13'h1bf9: q2 = 16'h48c2; // 0x37f2
	13'h1bfa: q2 = 16'hd3c2; // 0x37f4
	13'h1bfb: q2 = 16'hd3cb; // 0x37f6
	13'h1bfc: q2 = 16'h30a9; // 0x37f8
	13'h1bfd: q2 = 16'h0008; // 0x37fa
	13'h1bfe: q2 = 16'h5246; // 0x37fc
	13'h1bff: q2 = 16'h60ca; // 0x37fe
	13'h1c00: q2 = 16'h5247; // 0x3800
	13'h1c01: q2 = 16'h60be; // 0x3802
	13'h1c02: q2 = 16'h4246; // 0x3804
	13'h1c03: q2 = 16'hbc7c; // 0x3806
	13'h1c04: q2 = 16'h0004; // 0x3808
	13'h1c05: q2 = 16'h6c28; // 0x380a
	13'h1c06: q2 = 16'h3006; // 0x380c
	13'h1c07: q2 = 16'he340; // 0x380e
	13'h1c08: q2 = 16'h48c0; // 0x3810
	13'h1c09: q2 = 16'h2f00; // 0x3812
	13'h1c0a: q2 = 16'h3007; // 0x3814
	13'h1c0b: q2 = 16'he740; // 0x3816
	13'h1c0c: q2 = 16'h48c0; // 0x3818
	13'h1c0d: q2 = 16'h221f; // 0x381a
	13'h1c0e: q2 = 16'hd081; // 0x381c
	13'h1c0f: q2 = 16'hd08b; // 0x381e
	13'h1c10: q2 = 16'h2040; // 0x3820
	13'h1c11: q2 = 16'h3206; // 0x3822
	13'h1c12: q2 = 16'he341; // 0x3824
	13'h1c13: q2 = 16'h48c1; // 0x3826
	13'h1c14: q2 = 16'hd28e; // 0x3828
	13'h1c15: q2 = 16'h2241; // 0x382a
	13'h1c16: q2 = 16'h30a9; // 0x382c
	13'h1c17: q2 = 16'hff94; // 0x382e
	13'h1c18: q2 = 16'h5246; // 0x3830
	13'h1c19: q2 = 16'h60d2; // 0x3832
	13'h1c1a: q2 = 16'h3d7c; // 0x3834
	13'h1c1b: q2 = 16'h0002; // 0x3836
	13'h1c1c: q2 = 16'hffda; // 0x3838
	13'h1c1d: q2 = 16'h4247; // 0x383a
	13'h1c1e: q2 = 16'h2a7c; // 0x383c
	13'h1c1f: q2 = 16'h0000; // 0x383e
	13'h1c20: q2 = 16'hfe06; // 0x3840
	13'h1c21: q2 = 16'h287c; // 0x3842
	13'h1c22: q2 = 16'h0000; // 0x3844
	13'h1c23: q2 = 16'hfe16; // 0x3846
	13'h1c24: q2 = 16'hbe7c; // 0x3848
	13'h1c25: q2 = 16'h000f; // 0x384a
	13'h1c26: q2 = 16'h6c00; // 0x384c
	13'h1c27: q2 = 16'h00e6; // 0x384e
	13'h1c28: q2 = 16'h3007; // 0x3850
	13'h1c29: q2 = 16'he340; // 0x3852
	13'h1c2a: q2 = 16'h48c0; // 0x3854
	13'h1c2b: q2 = 16'hd08e; // 0x3856
	13'h1c2c: q2 = 16'h2040; // 0x3858
	13'h1c2d: q2 = 16'h4a68; // 0x385a
	13'h1c2e: q2 = 16'hffbc; // 0x385c
	13'h1c2f: q2 = 16'h6600; // 0x385e
	13'h1c30: q2 = 16'h00bc; // 0x3860
	13'h1c31: q2 = 16'h3007; // 0x3862
	13'h1c32: q2 = 16'he340; // 0x3864
	13'h1c33: q2 = 16'h48c0; // 0x3866
	13'h1c34: q2 = 16'hd08e; // 0x3868
	13'h1c35: q2 = 16'h2040; // 0x386a
	13'h1c36: q2 = 16'h5268; // 0x386c
	13'h1c37: q2 = 16'hff9e; // 0x386e
	13'h1c38: q2 = 16'h3007; // 0x3870
	13'h1c39: q2 = 16'he340; // 0x3872
	13'h1c3a: q2 = 16'h48c0; // 0x3874
	13'h1c3b: q2 = 16'hd08e; // 0x3876
	13'h1c3c: q2 = 16'h2040; // 0x3878
	13'h1c3d: q2 = 16'h0c68; // 0x387a
	13'h1c3e: q2 = 16'h000a; // 0x387c
	13'h1c3f: q2 = 16'hff9e; // 0x387e
	13'h1c40: q2 = 16'h6f16; // 0x3880
	13'h1c41: q2 = 16'h3007; // 0x3882
	13'h1c42: q2 = 16'he340; // 0x3884
	13'h1c43: q2 = 16'h48c0; // 0x3886
	13'h1c44: q2 = 16'hd08e; // 0x3888
	13'h1c45: q2 = 16'h2040; // 0x388a
	13'h1c46: q2 = 16'h4268; // 0x388c
	13'h1c47: q2 = 16'hff9e; // 0x388e
	13'h1c48: q2 = 16'h4a47; // 0x3890
	13'h1c49: q2 = 16'h6604; // 0x3892
	13'h1c4a: q2 = 16'h536e; // 0x3894
	13'h1c4b: q2 = 16'hff9c; // 0x3896
	13'h1c4c: q2 = 16'h3007; // 0x3898
	13'h1c4d: q2 = 16'he340; // 0x389a
	13'h1c4e: q2 = 16'h48c0; // 0x389c
	13'h1c4f: q2 = 16'hd08e; // 0x389e
	13'h1c50: q2 = 16'h2040; // 0x38a0
	13'h1c51: q2 = 16'h3207; // 0x38a2
	13'h1c52: q2 = 16'he341; // 0x38a4
	13'h1c53: q2 = 16'h48c1; // 0x38a6
	13'h1c54: q2 = 16'hd28e; // 0x38a8
	13'h1c55: q2 = 16'h2241; // 0x38aa
	13'h1c56: q2 = 16'h3229; // 0x38ac
	13'h1c57: q2 = 16'hff9e; // 0x38ae
	13'h1c58: q2 = 16'he341; // 0x38b0
	13'h1c59: q2 = 16'h48c1; // 0x38b2
	13'h1c5a: q2 = 16'hd2bc; // 0x38b4
	13'h1c5b: q2 = 16'h0000; // 0x38b6
	13'h1c5c: q2 = 16'hcab2; // 0x38b8
	13'h1c5d: q2 = 16'h2241; // 0x38ba
	13'h1c5e: q2 = 16'h3151; // 0x38bc
	13'h1c5f: q2 = 16'hffbc; // 0x38be
	13'h1c60: q2 = 16'h0c6e; // 0x38c0
	13'h1c61: q2 = 16'h0009; // 0x38c2
	13'h1c62: q2 = 16'hff9e; // 0x38c4
	13'h1c63: q2 = 16'h660c; // 0x38c6
	13'h1c64: q2 = 16'h2ebc; // 0x38c8
	13'h1c65: q2 = 16'h0000; // 0x38ca
	13'h1c66: q2 = 16'hc7bc; // 0x38cc
	13'h1c67: q2 = 16'h4eb9; // 0x38ce
	13'h1c68: q2 = 16'h0000; // 0x38d0
	13'h1c69: q2 = 16'h7dd8; // 0x38d2
	13'h1c6a: q2 = 16'h3e87; // 0x38d4
	13'h1c6b: q2 = 16'h0657; // 0x38d6
	13'h1c6c: q2 = 16'h0010; // 0x38d8
	13'h1c6d: q2 = 16'h3007; // 0x38da
	13'h1c6e: q2 = 16'he340; // 0x38dc
	13'h1c6f: q2 = 16'h48c0; // 0x38de
	13'h1c70: q2 = 16'hd08e; // 0x38e0
	13'h1c71: q2 = 16'h2040; // 0x38e2
	13'h1c72: q2 = 16'h3028; // 0x38e4
	13'h1c73: q2 = 16'hff9e; // 0x38e6
	13'h1c74: q2 = 16'he340; // 0x38e8
	13'h1c75: q2 = 16'h48c0; // 0x38ea
	13'h1c76: q2 = 16'hd0bc; // 0x38ec
	13'h1c77: q2 = 16'h0000; // 0x38ee
	13'h1c78: q2 = 16'hca9c; // 0x38f0
	13'h1c79: q2 = 16'h2040; // 0x38f2
	13'h1c7a: q2 = 16'h3f10; // 0x38f4
	13'h1c7b: q2 = 16'h1014; // 0x38f6
	13'h1c7c: q2 = 16'h4880; // 0x38f8
	13'h1c7d: q2 = 16'h3f00; // 0x38fa
	13'h1c7e: q2 = 16'h5357; // 0x38fc
	13'h1c7f: q2 = 16'h1015; // 0x38fe
	13'h1c80: q2 = 16'h4880; // 0x3900
	13'h1c81: q2 = 16'h3f00; // 0x3902
	13'h1c82: q2 = 16'hbe7c; // 0x3904
	13'h1c83: q2 = 16'h0003; // 0x3906
	13'h1c84: q2 = 16'h6c04; // 0x3908
	13'h1c85: q2 = 16'h700f; // 0x390a
	13'h1c86: q2 = 16'h6002; // 0x390c
	13'h1c87: q2 = 16'h700e; // 0x390e
	13'h1c88: q2 = 16'hd157; // 0x3910
	13'h1c89: q2 = 16'h4eb9; // 0x3912
	13'h1c8a: q2 = 16'h0000; // 0x3914
	13'h1c8b: q2 = 16'h3d18; // 0x3916
	13'h1c8c: q2 = 16'h5c4f; // 0x3918
	13'h1c8d: q2 = 16'h600e; // 0x391a
	13'h1c8e: q2 = 16'h3007; // 0x391c
	13'h1c8f: q2 = 16'he340; // 0x391e
	13'h1c90: q2 = 16'h48c0; // 0x3920
	13'h1c91: q2 = 16'hd08e; // 0x3922
	13'h1c92: q2 = 16'h2040; // 0x3924
	13'h1c93: q2 = 16'h5368; // 0x3926
	13'h1c94: q2 = 16'hffbc; // 0x3928
	13'h1c95: q2 = 16'h5247; // 0x392a
	13'h1c96: q2 = 16'h528d; // 0x392c
	13'h1c97: q2 = 16'h528c; // 0x392e
	13'h1c98: q2 = 16'h6000; // 0x3930
	13'h1c99: q2 = 16'hff16; // 0x3932
	13'h1c9a: q2 = 16'h4ab9; // 0x3934
	13'h1c9b: q2 = 16'h0001; // 0x3936
	13'h1c9c: q2 = 16'h7fc2; // 0x3938
	13'h1c9d: q2 = 16'h6720; // 0x393a
	13'h1c9e: q2 = 16'h4a6e; // 0x393c
	13'h1c9f: q2 = 16'hff9c; // 0x393e
	13'h1ca0: q2 = 16'h671e; // 0x3940
	13'h1ca1: q2 = 16'h4a79; // 0x3942
	13'h1ca2: q2 = 16'h0001; // 0x3944
	13'h1ca3: q2 = 16'h7f5e; // 0x3946
	13'h1ca4: q2 = 16'h6616; // 0x3948
	13'h1ca5: q2 = 16'h4a79; // 0x394a
	13'h1ca6: q2 = 16'h0001; // 0x394c
	13'h1ca7: q2 = 16'h7594; // 0x394e
	13'h1ca8: q2 = 16'h6708; // 0x3950
	13'h1ca9: q2 = 16'h4a79; // 0x3952
	13'h1caa: q2 = 16'h0001; // 0x3954
	13'h1cab: q2 = 16'h7fc6; // 0x3956
	13'h1cac: q2 = 16'h6606; // 0x3958
	13'h1cad: q2 = 16'h60d8; // 0x395a
	13'h1cae: q2 = 16'h6000; // 0x395c
	13'h1caf: q2 = 16'hfe26; // 0x395e
	13'h1cb0: q2 = 16'h4eb9; // 0x3960
	13'h1cb1: q2 = 16'h0000; // 0x3962
	13'h1cb2: q2 = 16'h0226; // 0x3964
	13'h1cb3: q2 = 16'h4eb9; // 0x3966
	13'h1cb4: q2 = 16'h0000; // 0x3968
	13'h1cb5: q2 = 16'h8ea8; // 0x396a
	13'h1cb6: q2 = 16'h4a9f; // 0x396c
	13'h1cb7: q2 = 16'h4cdf; // 0x396e
	13'h1cb8: q2 = 16'h38f0; // 0x3970
	13'h1cb9: q2 = 16'h4e5e; // 0x3972
	13'h1cba: q2 = 16'h4e75; // 0x3974
	13'h1cbb: q2 = 16'h4e56; // 0x3976
	13'h1cbc: q2 = 16'h0000; // 0x3978
	13'h1cbd: q2 = 16'h48e7; // 0x397a
	13'h1cbe: q2 = 16'h1f04; // 0x397c
	13'h1cbf: q2 = 16'h2e2e; // 0x397e
	13'h1cc0: q2 = 16'h0008; // 0x3980
	13'h1cc1: q2 = 16'h2a6e; // 0x3982
	13'h1cc2: q2 = 16'h000c; // 0x3984
	13'h1cc3: q2 = 16'h4215; // 0x3986
	13'h1cc4: q2 = 16'h2a3c; // 0x3988
	13'h1cc5: q2 = 16'h0000; // 0x398a
	13'h1cc6: q2 = 16'h0e10; // 0x398c
	13'h1cc7: q2 = 16'h7802; // 0x398e
	13'h1cc8: q2 = 16'h4a44; // 0x3990
	13'h1cc9: q2 = 16'h6d00; // 0x3992
	13'h1cca: q2 = 16'h008a; // 0x3994
	13'h1ccb: q2 = 16'hbe85; // 0x3996
	13'h1ccc: q2 = 16'h6f48; // 0x3998
	13'h1ccd: q2 = 16'h2f05; // 0x399a
	13'h1cce: q2 = 16'h2f07; // 0x399c
	13'h1ccf: q2 = 16'h4eb9; // 0x399e
	13'h1cd0: q2 = 16'h0000; // 0x39a0
	13'h1cd1: q2 = 16'h79ac; // 0x39a2
	13'h1cd2: q2 = 16'hbf8f; // 0x39a4
	13'h1cd3: q2 = 16'h2c00; // 0x39a6
	13'h1cd4: q2 = 16'hbcbc; // 0x39a8
	13'h1cd5: q2 = 16'h0000; // 0x39aa
	13'h1cd6: q2 = 16'h0009; // 0x39ac
	13'h1cd7: q2 = 16'h6c16; // 0x39ae
	13'h1cd8: q2 = 16'hb87c; // 0x39b0
	13'h1cd9: q2 = 16'h0002; // 0x39b2
	13'h1cda: q2 = 16'h6c10; // 0x39b4
	13'h1cdb: q2 = 16'h2ebc; // 0x39b6
	13'h1cdc: q2 = 16'h0000; // 0x39b8
	13'h1cdd: q2 = 16'hfe48; // 0x39ba
	13'h1cde: q2 = 16'h2f0d; // 0x39bc
	13'h1cdf: q2 = 16'h4eb9; // 0x39be
	13'h1ce0: q2 = 16'h0000; // 0x39c0
	13'h1ce1: q2 = 16'h0770; // 0x39c2
	13'h1ce2: q2 = 16'h4a9f; // 0x39c4
	13'h1ce3: q2 = 16'h2e8d; // 0x39c6
	13'h1ce4: q2 = 16'h2f06; // 0x39c8
	13'h1ce5: q2 = 16'h4eb9; // 0x39ca
	13'h1ce6: q2 = 16'h0000; // 0x39cc
	13'h1ce7: q2 = 16'h07c6; // 0x39ce
	13'h1ce8: q2 = 16'h4a9f; // 0x39d0
	13'h1ce9: q2 = 16'h2f05; // 0x39d2
	13'h1cea: q2 = 16'h2f06; // 0x39d4
	13'h1ceb: q2 = 16'h4eb9; // 0x39d6
	13'h1cec: q2 = 16'h0000; // 0x39d8
	13'h1ced: q2 = 16'h7a50; // 0x39da
	13'h1cee: q2 = 16'hbf8f; // 0x39dc
	13'h1cef: q2 = 16'h9e80; // 0x39de
	13'h1cf0: q2 = 16'h6010; // 0x39e0
	13'h1cf1: q2 = 16'h2ebc; // 0x39e2
	13'h1cf2: q2 = 16'h0000; // 0x39e4
	13'h1cf3: q2 = 16'hfe4a; // 0x39e6
	13'h1cf4: q2 = 16'h2f0d; // 0x39e8
	13'h1cf5: q2 = 16'h4eb9; // 0x39ea
	13'h1cf6: q2 = 16'h0000; // 0x39ec
	13'h1cf7: q2 = 16'h0770; // 0x39ee
	13'h1cf8: q2 = 16'h4a9f; // 0x39f0
	13'h1cf9: q2 = 16'h4a44; // 0x39f2
	13'h1cfa: q2 = 16'h6f10; // 0x39f4
	13'h1cfb: q2 = 16'h2ebc; // 0x39f6
	13'h1cfc: q2 = 16'h0000; // 0x39f8
	13'h1cfd: q2 = 16'hfe4d; // 0x39fa
	13'h1cfe: q2 = 16'h2f0d; // 0x39fc
	13'h1cff: q2 = 16'h4eb9; // 0x39fe
	13'h1d00: q2 = 16'h0000; // 0x3a00
	13'h1d01: q2 = 16'h0770; // 0x3a02
	13'h1d02: q2 = 16'h4a9f; // 0x3a04
	13'h1d03: q2 = 16'h2f39; // 0x3a06
	13'h1d04: q2 = 16'h0000; // 0x3a08
	13'h1d05: q2 = 16'hfe44; // 0x3a0a
	13'h1d06: q2 = 16'h2f05; // 0x3a0c
	13'h1d07: q2 = 16'h4eb9; // 0x3a0e
	13'h1d08: q2 = 16'h0000; // 0x3a10
	13'h1d09: q2 = 16'h79ac; // 0x3a12
	13'h1d0a: q2 = 16'hbf8f; // 0x3a14
	13'h1d0b: q2 = 16'h2a00; // 0x3a16
	13'h1d0c: q2 = 16'h5344; // 0x3a18
	13'h1d0d: q2 = 16'h6000; // 0x3a1a
	13'h1d0e: q2 = 16'hff74; // 0x3a1c
	13'h1d0f: q2 = 16'h4a9f; // 0x3a1e
	13'h1d10: q2 = 16'h4cdf; // 0x3a20
	13'h1d11: q2 = 16'h20f0; // 0x3a22
	13'h1d12: q2 = 16'h4e5e; // 0x3a24
	13'h1d13: q2 = 16'h4e75; // 0x3a26
	13'h1d14: q2 = 16'h207c; // 0x3a28
	13'h1d15: q2 = 16'h0001; // 0x3a2a
	13'h1d16: q2 = 16'h7a3e; // 0x3a2c
	13'h1d17: q2 = 16'h42a8; // 0x3a2e
	13'h1d18: q2 = 16'h000e; // 0x3a30
	13'h1d19: q2 = 16'h42a8; // 0x3a32
	13'h1d1a: q2 = 16'h0090; // 0x3a34
	13'h1d1b: q2 = 16'h4e75; // 0x3a36
	13'h1d1c: q2 = 16'h4e56; // 0x3a38
	13'h1d1d: q2 = 16'hfff6; // 0x3a3a
	13'h1d1e: q2 = 16'h2d7c; // 0x3a3c
	13'h1d1f: q2 = 16'h0001; // 0x3a3e
	13'h1d20: q2 = 16'h7a3e; // 0x3a40
	13'h1d21: q2 = 16'hfffc; // 0x3a42
	13'h1d22: q2 = 16'h6118; // 0x3a44
	13'h1d23: q2 = 16'h06ae; // 0x3a46
	13'h1d24: q2 = 16'h0000; // 0x3a48
	13'h1d25: q2 = 16'h0082; // 0x3a4a
	13'h1d26: q2 = 16'hfffc; // 0x3a4c
	13'h1d27: q2 = 16'h610e; // 0x3a4e
	13'h1d28: q2 = 16'h4e5e; // 0x3a50
	13'h1d29: q2 = 16'h5379; // 0x3a52
	13'h1d2a: q2 = 16'h0001; // 0x3a54
	13'h1d2b: q2 = 16'h7b9c; // 0x3a56
	13'h1d2c: q2 = 16'h6c00; // 0x3a58
	13'h1d2d: q2 = 16'hc5fc; // 0x3a5a
	13'h1d2e: q2 = 16'h4e75; // 0x3a5c
	13'h1d2f: q2 = 16'h206e; // 0x3a5e
	13'h1d30: q2 = 16'hfffc; // 0x3a60
	13'h1d31: q2 = 16'h4aa8; // 0x3a62
	13'h1d32: q2 = 16'h000e; // 0x3a64
	13'h1d33: q2 = 16'h67f4; // 0x3a66
	13'h1d34: q2 = 16'h2028; // 0x3a68
	13'h1d35: q2 = 16'h000a; // 0x3a6a
	13'h1d36: q2 = 16'hb0a8; // 0x3a6c
	13'h1d37: q2 = 16'h0004; // 0x3a6e
	13'h1d38: q2 = 16'h6f1a; // 0x3a70
	13'h1d39: q2 = 16'h206e; // 0x3a72
	13'h1d3a: q2 = 16'hfffc; // 0x3a74
	13'h1d3b: q2 = 16'h2028; // 0x3a76
	13'h1d3c: q2 = 16'h0000; // 0x3a78
	13'h1d3d: q2 = 16'hd1a8; // 0x3a7a
	13'h1d3e: q2 = 16'h0006; // 0x3a7c
	13'h1d3f: q2 = 16'h3028; // 0x3a7e
	13'h1d40: q2 = 16'h0004; // 0x3a80
	13'h1d41: q2 = 16'h4241; // 0x3a82
	13'h1d42: q2 = 16'hd141; // 0x3a84
	13'h1d43: q2 = 16'h3140; // 0x3a86
	13'h1d44: q2 = 16'h0004; // 0x3a88
	13'h1d45: q2 = 16'h4e75; // 0x3a8a
	13'h1d46: q2 = 16'h206e; // 0x3a8c
	13'h1d47: q2 = 16'hfffc; // 0x3a8e
	13'h1d48: q2 = 16'h2268; // 0x3a90
	13'h1d49: q2 = 16'h000e; // 0x3a92
	13'h1d4a: q2 = 16'h4240; // 0x3a94
	13'h1d4b: q2 = 16'h1019; // 0x3a96
	13'h1d4c: q2 = 16'h1d40; // 0x3a98
	13'h1d4d: q2 = 16'hfffb; // 0x3a9a
	13'h1d4e: q2 = 16'h2149; // 0x3a9c
	13'h1d4f: q2 = 16'h000e; // 0x3a9e
	13'h1d50: q2 = 16'h0880; // 0x3aa0
	13'h1d51: q2 = 16'h0007; // 0x3aa2
	13'h1d52: q2 = 16'he548; // 0x3aa4
	13'h1d53: q2 = 16'h247c; // 0x3aa6
	13'h1d54: q2 = 16'h0000; // 0x3aa8
	13'h1d55: q2 = 16'hfe50; // 0x3aaa
	13'h1d56: q2 = 16'hd4c0; // 0x3aac
	13'h1d57: q2 = 16'h2452; // 0x3aae
	13'h1d58: q2 = 16'h4e92; // 0x3ab0
	13'h1d59: q2 = 16'h082e; // 0x3ab2
	13'h1d5a: q2 = 16'h0007; // 0x3ab4
	13'h1d5b: q2 = 16'hfffb; // 0x3ab6
	13'h1d5c: q2 = 16'h67d2; // 0x3ab8
	13'h1d5d: q2 = 16'h206e; // 0x3aba
	13'h1d5e: q2 = 16'hfffc; // 0x3abc
	13'h1d5f: q2 = 16'h2268; // 0x3abe
	13'h1d60: q2 = 16'h000e; // 0x3ac0
	13'h1d61: q2 = 16'h4280; // 0x3ac2
	13'h1d62: q2 = 16'h3019; // 0x3ac4
	13'h1d63: q2 = 16'hd0a8; // 0x3ac6
	13'h1d64: q2 = 16'h000a; // 0x3ac8
	13'h1d65: q2 = 16'h640a; // 0x3aca
	13'h1d66: q2 = 16'h42a8; // 0x3acc
	13'h1d67: q2 = 16'h000a; // 0x3ace
	13'h1d68: q2 = 16'h42a8; // 0x3ad0
	13'h1d69: q2 = 16'h0004; // 0x3ad2
	13'h1d6a: q2 = 16'h60e8; // 0x3ad4
	13'h1d6b: q2 = 16'h2149; // 0x3ad6
	13'h1d6c: q2 = 16'h000e; // 0x3ad8
	13'h1d6d: q2 = 16'h2140; // 0x3ada
	13'h1d6e: q2 = 16'h000a; // 0x3adc
	13'h1d6f: q2 = 16'h6092; // 0x3ade
	13'h1d70: q2 = 16'h206e; // 0x3ae0
	13'h1d71: q2 = 16'hfffc; // 0x3ae2
	13'h1d72: q2 = 16'h2268; // 0x3ae4
	13'h1d73: q2 = 16'h000e; // 0x3ae6
	13'h1d74: q2 = 16'h1d59; // 0x3ae8
	13'h1d75: q2 = 16'hfffa; // 0x3aea
	13'h1d76: q2 = 16'h2149; // 0x3aec
	13'h1d77: q2 = 16'h000e; // 0x3aee
	13'h1d78: q2 = 16'hd1fc; // 0x3af0
	13'h1d79: q2 = 16'h0000; // 0x3af2
	13'h1d7a: q2 = 16'h001a; // 0x3af4
	13'h1d7b: q2 = 16'h2d48; // 0x3af6
	13'h1d7c: q2 = 16'hfff6; // 0x3af8
	13'h1d7d: q2 = 16'h082e; // 0x3afa
	13'h1d7e: q2 = 16'h0000; // 0x3afc
	13'h1d7f: q2 = 16'hfffa; // 0x3afe
	13'h1d80: q2 = 16'h6704; // 0x3b00
	13'h1d81: q2 = 16'h2057; // 0x3b02
	13'h1d82: q2 = 16'h4e90; // 0x3b04
	13'h1d83: q2 = 16'h06ae; // 0x3b06
	13'h1d84: q2 = 16'h0000; // 0x3b08
	13'h1d85: q2 = 16'h001a; // 0x3b0a
	13'h1d86: q2 = 16'hfff6; // 0x3b0c
	13'h1d87: q2 = 16'h102e; // 0x3b0e
	13'h1d88: q2 = 16'hfffa; // 0x3b10
	13'h1d89: q2 = 16'he208; // 0x3b12
	13'h1d8a: q2 = 16'h1d40; // 0x3b14
	13'h1d8b: q2 = 16'hfffa; // 0x3b16
	13'h1d8c: q2 = 16'h66e0; // 0x3b18
	13'h1d8d: q2 = 16'h588f; // 0x3b1a
	13'h1d8e: q2 = 16'h4e75; // 0x3b1c
	13'h1d8f: q2 = 16'h61c0; // 0x3b1e
	13'h1d90: q2 = 16'h3f3c; // 0x3b20
	13'h1d91: q2 = 16'hffff; // 0x3b22
	13'h1d92: q2 = 16'h2f2e; // 0x3b24
	13'h1d93: q2 = 16'hfff6; // 0x3b26
	13'h1d94: q2 = 16'h0697; // 0x3b28
	13'h1d95: q2 = 16'h0000; // 0x3b2a
	13'h1d96: q2 = 16'h000a; // 0x3b2c
	13'h1d97: q2 = 16'h3f3c; // 0x3b2e
	13'h1d98: q2 = 16'h0003; // 0x3b30
	13'h1d99: q2 = 16'h3f3c; // 0x3b32
	13'h1d9a: q2 = 16'h7530; // 0x3b34
	13'h1d9b: q2 = 16'h2f0f; // 0x3b36
	13'h1d9c: q2 = 16'h4eb9; // 0x3b38
	13'h1d9d: q2 = 16'h0000; // 0x3b3a
	13'h1d9e: q2 = 16'h7e06; // 0x3b3c
	13'h1d9f: q2 = 16'h4a40; // 0x3b3e
	13'h1da0: q2 = 16'h67fe; // 0x3b40
	13'h1da1: q2 = 16'hdffc; // 0x3b42
	13'h1da2: q2 = 16'h0000; // 0x3b44
	13'h1da3: q2 = 16'h000e; // 0x3b46
	13'h1da4: q2 = 16'h206e; // 0x3b48
	13'h1da5: q2 = 16'hfff6; // 0x3b4a
	13'h1da6: q2 = 16'h317c; // 0x3b4c
	13'h1da7: q2 = 16'h000c; // 0x3b4e
	13'h1da8: q2 = 16'h000c; // 0x3b50
	13'h1da9: q2 = 16'h3228; // 0x3b52
	13'h1daa: q2 = 16'h000a; // 0x3b54
	13'h1dab: q2 = 16'h227c; // 0x3b56
	13'h1dac: q2 = 16'h0000; // 0x3b58
	13'h1dad: q2 = 16'hca60; // 0x3b5a
	13'h1dae: q2 = 16'h3431; // 0x3b5c
	13'h1daf: q2 = 16'h1000; // 0x3b5e
	13'h1db0: q2 = 16'h247c; // 0x3b60
	13'h1db1: q2 = 16'h0001; // 0x3b62
	13'h1db2: q2 = 16'h7808; // 0x3b64
	13'h1db3: q2 = 16'h2588; // 0x3b66
	13'h1db4: q2 = 16'h2004; // 0x3b68
	13'h1db5: q2 = 16'h227c; // 0x3b6a
	13'h1db6: q2 = 16'h0000; // 0x3b6c
	13'h1db7: q2 = 16'hca7e; // 0x3b6e
	13'h1db8: q2 = 16'h3431; // 0x3b70
	13'h1db9: q2 = 16'h1000; // 0x3b72
	13'h1dba: q2 = 16'h35bc; // 0x3b74
	13'h1dbb: q2 = 16'h0001; // 0x3b76
	13'h1dbc: q2 = 16'h2000; // 0x3b78
	13'h1dbd: q2 = 16'h25bc; // 0x3b7a
	13'h1dbe: q2 = 16'h0040; // 0x3b7c
	13'h1dbf: q2 = 16'hffff; // 0x3b7e
	13'h1dc0: q2 = 16'h2004; // 0x3b80
	13'h1dc1: q2 = 16'h3431; // 0x3b82
	13'h1dc2: q2 = 16'h1002; // 0x3b84
	13'h1dc3: q2 = 16'h35bc; // 0x3b86
	13'h1dc4: q2 = 16'h0001; // 0x3b88
	13'h1dc5: q2 = 16'h2000; // 0x3b8a
	13'h1dc6: q2 = 16'h25bc; // 0x3b8c
	13'h1dc7: q2 = 16'h0020; // 0x3b8e
	13'h1dc8: q2 = 16'hffff; // 0x3b90
	13'h1dc9: q2 = 16'h2004; // 0x3b92
	13'h1dca: q2 = 16'h4e75; // 0x3b94
	13'h1dcb: q2 = 16'h206e; // 0x3b96
	13'h1dcc: q2 = 16'hfffc; // 0x3b98
	13'h1dcd: q2 = 16'h2028; // 0x3b9a
	13'h1dce: q2 = 16'h0016; // 0x3b9c
	13'h1dcf: q2 = 16'h2268; // 0x3b9e
	13'h1dd0: q2 = 16'h0012; // 0x3ba0
	13'h1dd1: q2 = 16'h4ed1; // 0x3ba2
	13'h1dd2: q2 = 16'h42a8; // 0x3ba4
	13'h1dd3: q2 = 16'h000e; // 0x3ba6
	13'h1dd4: q2 = 16'h584f; // 0x3ba8
	13'h1dd5: q2 = 16'h4e75; // 0x3baa
	13'h1dd6: q2 = 16'h206e; // 0x3bac
	13'h1dd7: q2 = 16'hfffc; // 0x3bae
	13'h1dd8: q2 = 16'h2268; // 0x3bb0
	13'h1dd9: q2 = 16'h000e; // 0x3bb2
	13'h1dda: q2 = 16'h5289; // 0x3bb4
	13'h1ddb: q2 = 16'h2159; // 0x3bb6
	13'h1ddc: q2 = 16'h0000; // 0x3bb8
	13'h1ddd: q2 = 16'h2149; // 0x3bba
	13'h1dde: q2 = 16'h000e; // 0x3bbc
	13'h1ddf: q2 = 16'h4e75; // 0x3bbe
	13'h1de0: q2 = 16'h720e; // 0x3bc0
	13'h1de1: q2 = 16'h6100; // 0x3bc2
	13'h1de2: q2 = 16'hff1c; // 0x3bc4
	13'h1de3: q2 = 16'h206e; // 0x3bc6
	13'h1de4: q2 = 16'hfffc; // 0x3bc8
	13'h1de5: q2 = 16'h226e; // 0x3bca
	13'h1de6: q2 = 16'hfff6; // 0x3bcc
	13'h1de7: q2 = 16'h2468; // 0x3bce
	13'h1de8: q2 = 16'h000e; // 0x3bd0
	13'h1de9: q2 = 16'h239a; // 0x3bd2
	13'h1dea: q2 = 16'h1000; // 0x3bd4
	13'h1deb: q2 = 16'h214a; // 0x3bd6
	13'h1dec: q2 = 16'h000e; // 0x3bd8
	13'h1ded: q2 = 16'h4e75; // 0x3bda
	13'h1dee: q2 = 16'h7212; // 0x3bdc
	13'h1def: q2 = 16'h60e2; // 0x3bde
	13'h1df0: q2 = 16'h7216; // 0x3be0
	13'h1df1: q2 = 16'h60de; // 0x3be2
	13'h1df2: q2 = 16'h6100; // 0x3be4
	13'h1df3: q2 = 16'hfefa; // 0x3be6
	13'h1df4: q2 = 16'h206e; // 0x3be8
	13'h1df5: q2 = 16'hfffc; // 0x3bea
	13'h1df6: q2 = 16'h226e; // 0x3bec
	13'h1df7: q2 = 16'hfff6; // 0x3bee
	13'h1df8: q2 = 16'h2468; // 0x3bf0
	13'h1df9: q2 = 16'h000e; // 0x3bf2
	13'h1dfa: q2 = 16'h235a; // 0x3bf4
	13'h1dfb: q2 = 16'h0000; // 0x3bf6
	13'h1dfc: q2 = 16'h670c; // 0x3bf8
	13'h1dfd: q2 = 16'h0069; // 0x3bfa
	13'h1dfe: q2 = 16'h0001; // 0x3bfc
	13'h1dff: q2 = 16'h000c; // 0x3bfe
	13'h1e00: q2 = 16'h214a; // 0x3c00
	13'h1e01: q2 = 16'h000e; // 0x3c02
	13'h1e02: q2 = 16'h4e75; // 0x3c04
	13'h1e03: q2 = 16'h0269; // 0x3c06
	13'h1e04: q2 = 16'hfffc; // 0x3c08
	13'h1e05: q2 = 16'h000c; // 0x3c0a
	13'h1e06: q2 = 16'h60f2; // 0x3c0c
	13'h1e07: q2 = 16'h6100; // 0x3c0e
	13'h1e08: q2 = 16'hfed0; // 0x3c10
	13'h1e09: q2 = 16'h610c; // 0x3c12
	13'h1e0a: q2 = 16'h206e; // 0x3c14
	13'h1e0b: q2 = 16'hfff6; // 0x3c16
	13'h1e0c: q2 = 16'h2268; // 0x3c18
	13'h1e0d: q2 = 16'h000e; // 0x3c1a
	13'h1e0e: q2 = 16'h6166; // 0x3c1c
	13'h1e0f: q2 = 16'h4e75; // 0x3c1e
	13'h1e10: q2 = 16'h206e; // 0x3c20
	13'h1e11: q2 = 16'hfff6; // 0x3c22
	13'h1e12: q2 = 16'h226e; // 0x3c24
	13'h1e13: q2 = 16'hfffc; // 0x3c26
	13'h1e14: q2 = 16'h2469; // 0x3c28
	13'h1e15: q2 = 16'h000e; // 0x3c2a
	13'h1e16: q2 = 16'h321a; // 0x3c2c
	13'h1e17: q2 = 16'h234a; // 0x3c2e
	13'h1e18: q2 = 16'h000e; // 0x3c30
	13'h1e19: q2 = 16'h3028; // 0x3c32
	13'h1e1a: q2 = 16'h000c; // 0x3c34
	13'h1e1b: q2 = 16'h0800; // 0x3c36
	13'h1e1c: q2 = 16'h0000; // 0x3c38
	13'h1e1d: q2 = 16'h6624; // 0x3c3a
	13'h1e1e: q2 = 16'h3141; // 0x3c3c
	13'h1e1f: q2 = 16'h0004; // 0x3c3e
	13'h1e20: q2 = 16'h4268; // 0x3c40
	13'h1e21: q2 = 16'h0006; // 0x3c42
	13'h1e22: q2 = 16'h247c; // 0x3c44
	13'h1e23: q2 = 16'h0000; // 0x3c46
	13'h1e24: q2 = 16'hbca4; // 0x3c48
	13'h1e25: q2 = 16'h227c; // 0x3c4a
	13'h1e26: q2 = 16'h0000; // 0x3c4c
	13'h1e27: q2 = 16'hca60; // 0x3c4e
	13'h1e28: q2 = 16'hd2e8; // 0x3c50
	13'h1e29: q2 = 16'h000a; // 0x3c52
	13'h1e2a: q2 = 16'h3251; // 0x3c54
	13'h1e2b: q2 = 16'hd3fc; // 0x3c56
	13'h1e2c: q2 = 16'h0001; // 0x3c58
	13'h1e2d: q2 = 16'h7808; // 0x3c5a
	13'h1e2e: q2 = 16'h228a; // 0x3c5c
	13'h1e2f: q2 = 16'h4e75; // 0x3c5e
	13'h1e30: q2 = 16'h0800; // 0x3c60
	13'h1e31: q2 = 16'h0001; // 0x3c62
	13'h1e32: q2 = 16'h6618; // 0x3c64
	13'h1e33: q2 = 16'hb268; // 0x3c66
	13'h1e34: q2 = 16'h0004; // 0x3c68
	13'h1e35: q2 = 16'h67f2; // 0x3c6a
	13'h1e36: q2 = 16'h247c; // 0x3c6c
	13'h1e37: q2 = 16'h0000; // 0x3c6e
	13'h1e38: q2 = 16'hbcb8; // 0x3c70
	13'h1e39: q2 = 16'h0068; // 0x3c72
	13'h1e3a: q2 = 16'h0002; // 0x3c74
	13'h1e3b: q2 = 16'h000c; // 0x3c76
	13'h1e3c: q2 = 16'h3141; // 0x3c78
	13'h1e3d: q2 = 16'h0008; // 0x3c7a
	13'h1e3e: q2 = 16'h60cc; // 0x3c7c
	13'h1e3f: q2 = 16'h3141; // 0x3c7e
	13'h1e40: q2 = 16'h0008; // 0x3c80
	13'h1e41: q2 = 16'h4e75; // 0x3c82
	13'h1e42: q2 = 16'h247c; // 0x3c84
	13'h1e43: q2 = 16'h0000; // 0x3c86
	13'h1e44: q2 = 16'hca60; // 0x3c88
	13'h1e45: q2 = 16'hd4e8; // 0x3c8a
	13'h1e46: q2 = 16'h000a; // 0x3c8c
	13'h1e47: q2 = 16'h3452; // 0x3c8e
	13'h1e48: q2 = 16'hd5fc; // 0x3c90
	13'h1e49: q2 = 16'h0001; // 0x3c92
	13'h1e4a: q2 = 16'h7808; // 0x3c94
	13'h1e4b: q2 = 16'hd4fc; // 0x3c96
	13'h1e4c: q2 = 16'h0038; // 0x3c98
	13'h1e4d: q2 = 16'h4cd9; // 0x3c9a
	13'h1e4e: q2 = 16'h0007; // 0x3c9c
	13'h1e4f: q2 = 16'h48e2; // 0x3c9e
	13'h1e50: q2 = 16'he000; // 0x3ca0
	13'h1e51: q2 = 16'h4e75; // 0x3ca2
	13'h1e52: q2 = 16'h206b; // 0x3ca4
	13'h1e53: q2 = 16'h0004; // 0x3ca6
	13'h1e54: q2 = 16'h4293; // 0x3ca8
	13'h1e55: q2 = 16'h1568; // 0x3caa
	13'h1e56: q2 = 16'h0004; // 0x3cac
	13'h1e57: q2 = 16'h0005; // 0x3cae
	13'h1e58: q2 = 16'h3028; // 0x3cb0
	13'h1e59: q2 = 16'h0004; // 0x3cb2
	13'h1e5a: q2 = 16'hef48; // 0x3cb4
	13'h1e5b: q2 = 16'h4e75; // 0x3cb6
	13'h1e5c: q2 = 16'h206b; // 0x3cb8
	13'h1e5d: q2 = 16'h0004; // 0x3cba
	13'h1e5e: q2 = 16'h3028; // 0x3cbc
	13'h1e5f: q2 = 16'h0004; // 0x3cbe
	13'h1e60: q2 = 16'hb068; // 0x3cc0
	13'h1e61: q2 = 16'h0008; // 0x3cc2
	13'h1e62: q2 = 16'h6e22; // 0x3cc4
	13'h1e63: q2 = 16'hc0e8; // 0x3cc6
	13'h1e64: q2 = 16'h0000; // 0x3cc8
	13'h1e65: q2 = 16'h4840; // 0x3cca
	13'h1e66: q2 = 16'hd068; // 0x3ccc
	13'h1e67: q2 = 16'h0004; // 0x3cce
	13'h1e68: q2 = 16'hb068; // 0x3cd0
	13'h1e69: q2 = 16'h0008; // 0x3cd2
	13'h1e6a: q2 = 16'h6d0c; // 0x3cd4
	13'h1e6b: q2 = 16'h3028; // 0x3cd6
	13'h1e6c: q2 = 16'h0008; // 0x3cd8
	13'h1e6d: q2 = 16'h0268; // 0x3cda
	13'h1e6e: q2 = 16'hfffd; // 0x3cdc
	13'h1e6f: q2 = 16'h000c; // 0x3cde
	13'h1e70: q2 = 16'h4293; // 0x3ce0
	13'h1e71: q2 = 16'h3140; // 0x3ce2
	13'h1e72: q2 = 16'h0004; // 0x3ce4
	13'h1e73: q2 = 16'h60c2; // 0x3ce6
	13'h1e74: q2 = 16'hc0e8; // 0x3ce8
	13'h1e75: q2 = 16'h0002; // 0x3cea
	13'h1e76: q2 = 16'h4840; // 0x3cec
	13'h1e77: q2 = 16'hb068; // 0x3cee
	13'h1e78: q2 = 16'h0008; // 0x3cf0
	13'h1e79: q2 = 16'h6eee; // 0x3cf2
	13'h1e7a: q2 = 16'h60e0; // 0x3cf4
	13'h1e7b: q2 = 16'h6100; // 0x3cf6
	13'h1e7c: q2 = 16'hfde8; // 0x3cf8
	13'h1e7d: q2 = 16'h206e; // 0x3cfa
	13'h1e7e: q2 = 16'hfff6; // 0x3cfc
	13'h1e7f: q2 = 16'h3268; // 0x3cfe
	13'h1e80: q2 = 16'h000a; // 0x3d00
	13'h1e81: q2 = 16'hd3fc; // 0x3d02
	13'h1e82: q2 = 16'h0001; // 0x3d04
	13'h1e83: q2 = 16'h7a00; // 0x3d06
	13'h1e84: q2 = 16'h3f11; // 0x3d08
	13'h1e85: q2 = 16'h4eb9; // 0x3d0a
	13'h1e86: q2 = 16'h0000; // 0x3d0c
	13'h1e87: q2 = 16'h824a; // 0x3d0e
	13'h1e88: q2 = 16'h548f; // 0x3d10
	13'h1e89: q2 = 16'h4e75; // 0x3d12
	13'h1e8a: q2 = 16'h6100; // 0x3d14
	13'h1e8b: q2 = 16'hfdca; // 0x3d16
	13'h1e8c: q2 = 16'h6100; // 0x3d18
	13'h1e8d: q2 = 16'hff06; // 0x3d1a
	13'h1e8e: q2 = 16'h206e; // 0x3d1c
	13'h1e8f: q2 = 16'hfff6; // 0x3d1e
	13'h1e90: q2 = 16'h2268; // 0x3d20
	13'h1e91: q2 = 16'h0012; // 0x3d22
	13'h1e92: q2 = 16'h6100; // 0x3d24
	13'h1e93: q2 = 16'hff5e; // 0x3d26
	13'h1e94: q2 = 16'h4e75; // 0x3d28
	13'h1e95: q2 = 16'h6100; // 0x3d2a
	13'h1e96: q2 = 16'hfdb4; // 0x3d2c
	13'h1e97: q2 = 16'h206e; // 0x3d2e
	13'h1e98: q2 = 16'hfff6; // 0x3d30
	13'h1e99: q2 = 16'h2268; // 0x3d32
	13'h1e9a: q2 = 16'h0016; // 0x3d34
	13'h1e9b: q2 = 16'h6100; // 0x3d36
	13'h1e9c: q2 = 16'hff4c; // 0x3d38
	13'h1e9d: q2 = 16'h4e75; // 0x3d3a
	13'h1e9e: q2 = 16'h6100; // 0x3d3c
	13'h1e9f: q2 = 16'hfda2; // 0x3d3e
	13'h1ea0: q2 = 16'h6100; // 0x3d40
	13'h1ea1: q2 = 16'hfede; // 0x3d42
	13'h1ea2: q2 = 16'h4e75; // 0x3d44
	13'h1ea3: q2 = 16'h206e; // 0x3d46
	13'h1ea4: q2 = 16'hfffc; // 0x3d48
	13'h1ea5: q2 = 16'h52a8; // 0x3d4a
	13'h1ea6: q2 = 16'h000e; // 0x3d4c
	13'h1ea7: q2 = 16'h4e75; // 0x3d4e
	13'h1ea8: q2 = 16'h206e; // 0x3d50
	13'h1ea9: q2 = 16'hfffc; // 0x3d52
	13'h1eaa: q2 = 16'h217c; // 0x3d54
	13'h1eab: q2 = 16'h0000; // 0x3d56
	13'h1eac: q2 = 16'hbd6c; // 0x3d58
	13'h1ead: q2 = 16'h0012; // 0x3d5a
	13'h1eae: q2 = 16'h2268; // 0x3d5c
	13'h1eaf: q2 = 16'h000e; // 0x3d5e
	13'h1eb0: q2 = 16'h5289; // 0x3d60
	13'h1eb1: q2 = 16'h2159; // 0x3d62
	13'h1eb2: q2 = 16'h000e; // 0x3d64
	13'h1eb3: q2 = 16'h2149; // 0x3d66
	13'h1eb4: q2 = 16'h0016; // 0x3d68
	13'h1eb5: q2 = 16'h4e75; // 0x3d6a
	13'h1eb6: q2 = 16'h206e; // 0x3d6c
	13'h1eb7: q2 = 16'hfffc; // 0x3d6e
	13'h1eb8: q2 = 16'h2140; // 0x3d70
	13'h1eb9: q2 = 16'h000e; // 0x3d72
	13'h1eba: q2 = 16'h217c; // 0x3d74
	13'h1ebb: q2 = 16'h0000; // 0x3d76
	13'h1ebc: q2 = 16'hbba4; // 0x3d78
	13'h1ebd: q2 = 16'h0012; // 0x3d7a
	13'h1ebe: q2 = 16'h4e75; // 0x3d7c
	13'h1ebf: q2 = 16'h206e; // 0x3d7e
	13'h1ec0: q2 = 16'hfffc; // 0x3d80
	13'h1ec1: q2 = 16'h2268; // 0x3d82
	13'h1ec2: q2 = 16'h000e; // 0x3d84
	13'h1ec3: q2 = 16'h5289; // 0x3d86
	13'h1ec4: q2 = 16'h2f19; // 0x3d88
	13'h1ec5: q2 = 16'h2149; // 0x3d8a
	13'h1ec6: q2 = 16'h000e; // 0x3d8c
	13'h1ec7: q2 = 16'h4eb9; // 0x3d8e
	13'h1ec8: q2 = 16'h0000; // 0x3d90
	13'h1ec9: q2 = 16'h7e06; // 0x3d92
	13'h1eca: q2 = 16'h588f; // 0x3d94
	13'h1ecb: q2 = 16'h4e75; // 0x3d96
	13'h1ecc: q2 = 16'h206e; // 0x3d98
	13'h1ecd: q2 = 16'hfffc; // 0x3d9a
	13'h1ece: q2 = 16'h52a8; // 0x3d9c
	13'h1ecf: q2 = 16'h000e; // 0x3d9e
	13'h1ed0: q2 = 16'h33fc; // 0x3da0
	13'h1ed1: q2 = 16'h0000; // 0x3da2
	13'h1ed2: q2 = 16'h0001; // 0x3da4
	13'h1ed3: q2 = 16'h86a8; // 0x3da6
	13'h1ed4: q2 = 16'h4e75; // 0x3da8
	13'h1ed5: q2 = 16'h4e56; // 0x3daa
	13'h1ed6: q2 = 16'h0000; // 0x3dac
	13'h1ed7: q2 = 16'h48e7; // 0x3dae
	13'h1ed8: q2 = 16'h0f1c; // 0x3db0
	13'h1ed9: q2 = 16'h2a7c; // 0x3db2
	13'h1eda: q2 = 16'h0001; // 0x3db4
	13'h1edb: q2 = 16'h7f64; // 0x3db6
	13'h1edc: q2 = 16'h287c; // 0x3db8
	13'h1edd: q2 = 16'h0001; // 0x3dba
	13'h1ede: q2 = 16'h7ba8; // 0x3dbc
	13'h1edf: q2 = 16'h267c; // 0x3dbe
	13'h1ee0: q2 = 16'h0001; // 0x3dc0
	13'h1ee1: q2 = 16'h7efe; // 0x3dc2
	13'h1ee2: q2 = 16'h302e; // 0x3dc4
	13'h1ee3: q2 = 16'h0008; // 0x3dc6
	13'h1ee4: q2 = 16'hc1fc; // 0x3dc8
	13'h1ee5: q2 = 16'h0026; // 0x3dca
	13'h1ee6: q2 = 16'hd0bc; // 0x3dcc
	13'h1ee7: q2 = 16'h0001; // 0x3dce
	13'h1ee8: q2 = 16'h862c; // 0x3dd0
	13'h1ee9: q2 = 16'h2040; // 0x3dd2
	13'h1eea: q2 = 16'h2a10; // 0x3dd4
	13'h1eeb: q2 = 16'hbaad; // 0x3dd6
	13'h1eec: q2 = 16'h0038; // 0x3dd8
	13'h1eed: q2 = 16'h6f00; // 0x3dda
	13'h1eee: q2 = 16'h00fa; // 0x3ddc
	13'h1eef: q2 = 16'h7e0e; // 0x3dde
	13'h1ef0: q2 = 16'h4a47; // 0x3de0
	13'h1ef1: q2 = 16'h6716; // 0x3de2
	13'h1ef2: q2 = 16'h3007; // 0x3de4
	13'h1ef3: q2 = 16'h5340; // 0x3de6
	13'h1ef4: q2 = 16'he540; // 0x3de8
	13'h1ef5: q2 = 16'h48c0; // 0x3dea
	13'h1ef6: q2 = 16'hd08d; // 0x3dec
	13'h1ef7: q2 = 16'h2040; // 0x3dee
	13'h1ef8: q2 = 16'h2010; // 0x3df0
	13'h1ef9: q2 = 16'hb085; // 0x3df2
	13'h1efa: q2 = 16'h6c04; // 0x3df4
	13'h1efb: q2 = 16'h5347; // 0x3df6
	13'h1efc: q2 = 16'h60e6; // 0x3df8
	13'h1efd: q2 = 16'h7c29; // 0x3dfa
	13'h1efe: q2 = 16'h3007; // 0x3dfc
	13'h1eff: q2 = 16'hc1fc; // 0x3dfe
	13'h1f00: q2 = 16'h0003; // 0x3e00
	13'h1f01: q2 = 16'hb046; // 0x3e02
	13'h1f02: q2 = 16'h6e1c; // 0x3e04
	13'h1f03: q2 = 16'h3206; // 0x3e06
	13'h1f04: q2 = 16'h48c1; // 0x3e08
	13'h1f05: q2 = 16'h200c; // 0x3e0a
	13'h1f06: q2 = 16'hd081; // 0x3e0c
	13'h1f07: q2 = 16'h2040; // 0x3e0e
	13'h1f08: q2 = 16'h3406; // 0x3e10
	13'h1f09: q2 = 16'h48c2; // 0x3e12
	13'h1f0a: q2 = 16'h220c; // 0x3e14
	13'h1f0b: q2 = 16'hd282; // 0x3e16
	13'h1f0c: q2 = 16'h2241; // 0x3e18
	13'h1f0d: q2 = 16'h1151; // 0x3e1a
	13'h1f0e: q2 = 16'h0003; // 0x3e1c
	13'h1f0f: q2 = 16'h5346; // 0x3e1e
	13'h1f10: q2 = 16'h60da; // 0x3e20
	13'h1f11: q2 = 16'h7c0d; // 0x3e22
	13'h1f12: q2 = 16'hbc47; // 0x3e24
	13'h1f13: q2 = 16'h6d34; // 0x3e26
	13'h1f14: q2 = 16'h3006; // 0x3e28
	13'h1f15: q2 = 16'he540; // 0x3e2a
	13'h1f16: q2 = 16'h48c0; // 0x3e2c
	13'h1f17: q2 = 16'hd08d; // 0x3e2e
	13'h1f18: q2 = 16'h2040; // 0x3e30
	13'h1f19: q2 = 16'h3206; // 0x3e32
	13'h1f1a: q2 = 16'he541; // 0x3e34
	13'h1f1b: q2 = 16'h48c1; // 0x3e36
	13'h1f1c: q2 = 16'hd28d; // 0x3e38
	13'h1f1d: q2 = 16'h2241; // 0x3e3a
	13'h1f1e: q2 = 16'h2350; // 0x3e3c
	13'h1f1f: q2 = 16'h0004; // 0x3e3e
	13'h1f20: q2 = 16'h3006; // 0x3e40
	13'h1f21: q2 = 16'he340; // 0x3e42
	13'h1f22: q2 = 16'h48c0; // 0x3e44
	13'h1f23: q2 = 16'hd08b; // 0x3e46
	13'h1f24: q2 = 16'h2040; // 0x3e48
	13'h1f25: q2 = 16'h3206; // 0x3e4a
	13'h1f26: q2 = 16'he341; // 0x3e4c
	13'h1f27: q2 = 16'h48c1; // 0x3e4e
	13'h1f28: q2 = 16'hd28b; // 0x3e50
	13'h1f29: q2 = 16'h2241; // 0x3e52
	13'h1f2a: q2 = 16'h3151; // 0x3e54
	13'h1f2b: q2 = 16'h0002; // 0x3e56
	13'h1f2c: q2 = 16'h5346; // 0x3e58
	13'h1f2d: q2 = 16'h60c8; // 0x3e5a
	13'h1f2e: q2 = 16'h3007; // 0x3e5c
	13'h1f2f: q2 = 16'he540; // 0x3e5e
	13'h1f30: q2 = 16'h48c0; // 0x3e60
	13'h1f31: q2 = 16'hd08d; // 0x3e62
	13'h1f32: q2 = 16'h2040; // 0x3e64
	13'h1f33: q2 = 16'h2085; // 0x3e66
	13'h1f34: q2 = 16'h3007; // 0x3e68
	13'h1f35: q2 = 16'he340; // 0x3e6a
	13'h1f36: q2 = 16'h48c0; // 0x3e6c
	13'h1f37: q2 = 16'hd08b; // 0x3e6e
	13'h1f38: q2 = 16'h2040; // 0x3e70
	13'h1f39: q2 = 16'h322e; // 0x3e72
	13'h1f3a: q2 = 16'h0008; // 0x3e74
	13'h1f3b: q2 = 16'hc3fc; // 0x3e76
	13'h1f3c: q2 = 16'h0026; // 0x3e78
	13'h1f3d: q2 = 16'hd2bc; // 0x3e7a
	13'h1f3e: q2 = 16'h0001; // 0x3e7c
	13'h1f3f: q2 = 16'h8628; // 0x3e7e
	13'h1f40: q2 = 16'h2241; // 0x3e80
	13'h1f41: q2 = 16'h3091; // 0x3e82
	13'h1f42: q2 = 16'h3007; // 0x3e84
	13'h1f43: q2 = 16'hc1fc; // 0x3e86
	13'h1f44: q2 = 16'h0003; // 0x3e88
	13'h1f45: q2 = 16'h48c0; // 0x3e8a
	13'h1f46: q2 = 16'hd9c0; // 0x3e8c
	13'h1f47: q2 = 16'h18bc; // 0x3e8e
	13'h1f48: q2 = 16'h0047; // 0x3e90
	13'h1f49: q2 = 16'h197c; // 0x3e92
	13'h1f4a: q2 = 16'h0043; // 0x3e94
	13'h1f4b: q2 = 16'h0001; // 0x3e96
	13'h1f4c: q2 = 16'h197c; // 0x3e98
	13'h1f4d: q2 = 16'h0043; // 0x3e9a
	13'h1f4e: q2 = 16'h0002; // 0x3e9c
	13'h1f4f: q2 = 16'h302e; // 0x3e9e
	13'h1f50: q2 = 16'h0008; // 0x3ea0
	13'h1f51: q2 = 16'hc1fc; // 0x3ea2
	13'h1f52: q2 = 16'h0026; // 0x3ea4
	13'h1f53: q2 = 16'hd0bc; // 0x3ea6
	13'h1f54: q2 = 16'h0001; // 0x3ea8
	13'h1f55: q2 = 16'h8646; // 0x3eaa
	13'h1f56: q2 = 16'h2040; // 0x3eac
	13'h1f57: q2 = 16'h3207; // 0x3eae
	13'h1f58: q2 = 16'h5241; // 0x3eb0
	13'h1f59: q2 = 16'h3081; // 0x3eb2
	13'h1f5a: q2 = 16'h4a47; // 0x3eb4
	13'h1f5b: q2 = 16'h661e; // 0x3eb6
	13'h1f5c: q2 = 16'h302e; // 0x3eb8
	13'h1f5d: q2 = 16'h0008; // 0x3eba
	13'h1f5e: q2 = 16'hc1fc; // 0x3ebc
	13'h1f5f: q2 = 16'h0026; // 0x3ebe
	13'h1f60: q2 = 16'hd0bc; // 0x3ec0
	13'h1f61: q2 = 16'h0001; // 0x3ec2
	13'h1f62: q2 = 16'h8630; // 0x3ec4
	13'h1f63: q2 = 16'h2e80; // 0x3ec6
	13'h1f64: q2 = 16'h2f3c; // 0x3ec8
	13'h1f65: q2 = 16'h0001; // 0x3eca
	13'h1f66: q2 = 16'h860e; // 0x3ecc
	13'h1f67: q2 = 16'h4eb9; // 0x3ece
	13'h1f68: q2 = 16'h0000; // 0x3ed0
	13'h1f69: q2 = 16'h0750; // 0x3ed2
	13'h1f6a: q2 = 16'h4a9f; // 0x3ed4
	13'h1f6b: q2 = 16'h4a9f; // 0x3ed6
	13'h1f6c: q2 = 16'h4cdf; // 0x3ed8
	13'h1f6d: q2 = 16'h38e0; // 0x3eda
	13'h1f6e: q2 = 16'h4e5e; // 0x3edc
	13'h1f6f: q2 = 16'h4e75; // 0x3ede
	13'h1f70: q2 = 16'h4e56; // 0x3ee0
	13'h1f71: q2 = 16'h0000; // 0x3ee2
	13'h1f72: q2 = 16'h48e7; // 0x3ee4
	13'h1f73: q2 = 16'h010c; // 0x3ee6
	13'h1f74: q2 = 16'h2a6e; // 0x3ee8
	13'h1f75: q2 = 16'h0008; // 0x3eea
	13'h1f76: q2 = 16'h286e; // 0x3eec
	13'h1f77: q2 = 16'h000c; // 0x3eee
	13'h1f78: q2 = 16'h3015; // 0x3ef0
	13'h1f79: q2 = 16'hee40; // 0x3ef2
	13'h1f7a: q2 = 16'h3a80; // 0x3ef4
	13'h1f7b: q2 = 16'h3015; // 0x3ef6
	13'h1f7c: q2 = 16'h5340; // 0x3ef8
	13'h1f7d: q2 = 16'h3a80; // 0x3efa
	13'h1f7e: q2 = 16'h3015; // 0x3efc
	13'h1f7f: q2 = 16'hc07c; // 0x3efe
	13'h1f80: q2 = 16'hfff8; // 0x3f00
	13'h1f81: q2 = 16'h3a80; // 0x3f02
	13'h1f82: q2 = 16'h3015; // 0x3f04
	13'h1f83: q2 = 16'hef40; // 0x3f06
	13'h1f84: q2 = 16'h3a80; // 0x3f08
	13'h1f85: q2 = 16'h3014; // 0x3f0a
	13'h1f86: q2 = 16'hee40; // 0x3f0c
	13'h1f87: q2 = 16'hc07c; // 0x3f0e
	13'h1f88: q2 = 16'hfff8; // 0x3f10
	13'h1f89: q2 = 16'hef40; // 0x3f12
	13'h1f8a: q2 = 16'h3880; // 0x3f14
	13'h1f8b: q2 = 16'h4a9f; // 0x3f16
	13'h1f8c: q2 = 16'h4cdf; // 0x3f18
	13'h1f8d: q2 = 16'h3000; // 0x3f1a
	13'h1f8e: q2 = 16'h4e5e; // 0x3f1c
	13'h1f8f: q2 = 16'h4e75; // 0x3f1e
	13'h1f90: q2 = 16'h2021; // 0x3f20
	13'h1f91: q2 = 16'h2223; // 0x3f22
	13'h1f92: q2 = 16'h2425; // 0x3f24
	13'h1f93: q2 = 16'h2627; // 0x3f26
	13'h1f94: q2 = 16'h2829; // 0x3f28
	13'h1f95: q2 = 16'h2a2b; // 0x3f2a
	13'h1f96: q2 = 16'h2c2d; // 0x3f2c
	13'h1f97: q2 = 16'h2e2f; // 0x3f2e
	13'h1f98: q2 = 16'h3031; // 0x3f30
	13'h1f99: q2 = 16'h3233; // 0x3f32
	13'h1f9a: q2 = 16'h3435; // 0x3f34
	13'h1f9b: q2 = 16'h3637; // 0x3f36
	13'h1f9c: q2 = 16'h3839; // 0x3f38
	13'h1f9d: q2 = 16'h3a3b; // 0x3f3a
	13'h1f9e: q2 = 16'h3c3d; // 0x3f3c
	13'h1f9f: q2 = 16'h3e3f; // 0x3f3e
	13'h1fa0: q2 = 16'h4041; // 0x3f40
	13'h1fa1: q2 = 16'h4243; // 0x3f42
	13'h1fa2: q2 = 16'h4445; // 0x3f44
	13'h1fa3: q2 = 16'h4647; // 0x3f46
	13'h1fa4: q2 = 16'h4849; // 0x3f48
	13'h1fa5: q2 = 16'h4a4b; // 0x3f4a
	13'h1fa6: q2 = 16'h4c4d; // 0x3f4c
	13'h1fa7: q2 = 16'h4e4f; // 0x3f4e
	13'h1fa8: q2 = 16'h5051; // 0x3f50
	13'h1fa9: q2 = 16'h5253; // 0x3f52
	13'h1faa: q2 = 16'h5455; // 0x3f54
	13'h1fab: q2 = 16'h5657; // 0x3f56
	13'h1fac: q2 = 16'h5859; // 0x3f58
	13'h1fad: q2 = 16'h5a5b; // 0x3f5a
	13'h1fae: q2 = 16'h5c5d; // 0x3f5c
	13'h1faf: q2 = 16'h5e5f; // 0x3f5e
	13'h1fb0: q2 = 16'h6061; // 0x3f60
	13'h1fb1: q2 = 16'h6263; // 0x3f62
	13'h1fb2: q2 = 16'h6465; // 0x3f64
	13'h1fb3: q2 = 16'h6667; // 0x3f66
	13'h1fb4: q2 = 16'h6869; // 0x3f68
	13'h1fb5: q2 = 16'h6a6b; // 0x3f6a
	13'h1fb6: q2 = 16'h6c6d; // 0x3f6c
	13'h1fb7: q2 = 16'h6e6f; // 0x3f6e
	13'h1fb8: q2 = 16'h7071; // 0x3f70
	13'h1fb9: q2 = 16'h7273; // 0x3f72
	13'h1fba: q2 = 16'h7475; // 0x3f74
	13'h1fbb: q2 = 16'h7677; // 0x3f76
	13'h1fbc: q2 = 16'h7879; // 0x3f78
	13'h1fbd: q2 = 16'h7a7b; // 0x3f7a
	13'h1fbe: q2 = 16'h7c7d; // 0x3f7c
	13'h1fbf: q2 = 16'h7e7f; // 0x3f7e
	13'h1fc0: q2 = 16'h8081; // 0x3f80
	13'h1fc1: q2 = 16'h8283; // 0x3f82
	13'h1fc2: q2 = 16'h8485; // 0x3f84
	13'h1fc3: q2 = 16'h8687; // 0x3f86
	13'h1fc4: q2 = 16'h8889; // 0x3f88
	13'h1fc5: q2 = 16'h8a8b; // 0x3f8a
	13'h1fc6: q2 = 16'h8c8d; // 0x3f8c
	13'h1fc7: q2 = 16'h8e8f; // 0x3f8e
	13'h1fc8: q2 = 16'h9091; // 0x3f90
	13'h1fc9: q2 = 16'h9293; // 0x3f92
	13'h1fca: q2 = 16'h9495; // 0x3f94
	13'h1fcb: q2 = 16'h9697; // 0x3f96
	13'h1fcc: q2 = 16'h9899; // 0x3f98
	13'h1fcd: q2 = 16'h9a9b; // 0x3f9a
	13'h1fce: q2 = 16'h9c9d; // 0x3f9c
	13'h1fcf: q2 = 16'h9e9f; // 0x3f9e
	13'h1fd0: q2 = 16'ha0a1; // 0x3fa0
	13'h1fd1: q2 = 16'ha2a3; // 0x3fa2
	13'h1fd2: q2 = 16'ha4a5; // 0x3fa4
	13'h1fd3: q2 = 16'ha6a7; // 0x3fa6
	13'h1fd4: q2 = 16'ha8a9; // 0x3fa8
	13'h1fd5: q2 = 16'haaab; // 0x3faa
	13'h1fd6: q2 = 16'hacad; // 0x3fac
	13'h1fd7: q2 = 16'haeaf; // 0x3fae
	13'h1fd8: q2 = 16'hb0b1; // 0x3fb0
	13'h1fd9: q2 = 16'hb2b3; // 0x3fb2
	13'h1fda: q2 = 16'hb4b5; // 0x3fb4
	13'h1fdb: q2 = 16'hb6b7; // 0x3fb6
	13'h1fdc: q2 = 16'hb8b9; // 0x3fb8
	13'h1fdd: q2 = 16'hbabb; // 0x3fba
	13'h1fde: q2 = 16'hbcbd; // 0x3fbc
	13'h1fdf: q2 = 16'hbebf; // 0x3fbe
	13'h1fe0: q2 = 16'hc0c1; // 0x3fc0
	13'h1fe1: q2 = 16'hc2c3; // 0x3fc2
	13'h1fe2: q2 = 16'hc4c5; // 0x3fc4
	13'h1fe3: q2 = 16'hc6c7; // 0x3fc6
	13'h1fe4: q2 = 16'hc8c9; // 0x3fc8
	13'h1fe5: q2 = 16'hcacb; // 0x3fca
	13'h1fe6: q2 = 16'hcccd; // 0x3fcc
	13'h1fe7: q2 = 16'hcecf; // 0x3fce
	13'h1fe8: q2 = 16'hd0d1; // 0x3fd0
	13'h1fe9: q2 = 16'hd2d3; // 0x3fd2
	13'h1fea: q2 = 16'hd4d5; // 0x3fd4
	13'h1feb: q2 = 16'hd6d7; // 0x3fd6
	13'h1fec: q2 = 16'hd8d9; // 0x3fd8
	13'h1fed: q2 = 16'hdadb; // 0x3fda
	13'h1fee: q2 = 16'hdcdd; // 0x3fdc
	13'h1fef: q2 = 16'hdedf; // 0x3fde
	13'h1ff0: q2 = 16'he0e1; // 0x3fe0
	13'h1ff1: q2 = 16'he2e3; // 0x3fe2
	13'h1ff2: q2 = 16'he4e5; // 0x3fe4
	13'h1ff3: q2 = 16'he6e7; // 0x3fe6
	13'h1ff4: q2 = 16'he8e9; // 0x3fe8
	13'h1ff5: q2 = 16'heaeb; // 0x3fea
	13'h1ff6: q2 = 16'heced; // 0x3fec
	13'h1ff7: q2 = 16'heeef; // 0x3fee
	13'h1ff8: q2 = 16'hf0f1; // 0x3ff0
	13'h1ff9: q2 = 16'hf2f3; // 0x3ff2
	13'h1ffa: q2 = 16'hf4f5; // 0x3ff4
	13'h1ffb: q2 = 16'hf6f7; // 0x3ff6
	13'h1ffc: q2 = 16'hf8f9; // 0x3ff8
	13'h1ffd: q2 = 16'hfafb; // 0x3ffa
	13'h1ffe: q2 = 16'hfcfd; // 0x3ffc
	13'h1fff: q2 = 16'hfeff; // 0x3ffe
  endcase

  always @(posedge clk)
    case (a)
	// foodfight code 136020-208.9f, 136020-307.8f
	13'h0000: q3 = 16'h0001; // 0x0000
	13'h0001: q3 = 16'h0203; // 0x0002
	13'h0002: q3 = 16'h0405; // 0x0004
	13'h0003: q3 = 16'h0607; // 0x0006
	13'h0004: q3 = 16'h0809; // 0x0008
	13'h0005: q3 = 16'h0a0b; // 0x000a
	13'h0006: q3 = 16'h0c0d; // 0x000c
	13'h0007: q3 = 16'h0e0f; // 0x000e
	13'h0008: q3 = 16'h1011; // 0x0010
	13'h0009: q3 = 16'h1213; // 0x0012
	13'h000a: q3 = 16'h1415; // 0x0014
	13'h000b: q3 = 16'h1617; // 0x0016
	13'h000c: q3 = 16'h1819; // 0x0018
	13'h000d: q3 = 16'h1a1b; // 0x001a
	13'h000e: q3 = 16'h1c1d; // 0x001c
	13'h000f: q3 = 16'h1e1f; // 0x001e
	13'h0010: q3 = 16'h2021; // 0x0020
	13'h0011: q3 = 16'h2223; // 0x0022
	13'h0012: q3 = 16'h2425; // 0x0024
	13'h0013: q3 = 16'h2627; // 0x0026
	13'h0014: q3 = 16'h2829; // 0x0028
	13'h0015: q3 = 16'h2a2b; // 0x002a
	13'h0016: q3 = 16'h2c2d; // 0x002c
	13'h0017: q3 = 16'h2e2f; // 0x002e
	13'h0018: q3 = 16'h3031; // 0x0030
	13'h0019: q3 = 16'h3233; // 0x0032
	13'h001a: q3 = 16'h3435; // 0x0034
	13'h001b: q3 = 16'h3637; // 0x0036
	13'h001c: q3 = 16'h3839; // 0x0038
	13'h001d: q3 = 16'h3a3b; // 0x003a
	13'h001e: q3 = 16'h3c3d; // 0x003c
	13'h001f: q3 = 16'h3e3f; // 0x003e
	13'h0020: q3 = 16'h4041; // 0x0040
	13'h0021: q3 = 16'h4243; // 0x0042
	13'h0022: q3 = 16'h4445; // 0x0044
	13'h0023: q3 = 16'h4647; // 0x0046
	13'h0024: q3 = 16'h4849; // 0x0048
	13'h0025: q3 = 16'h4a4b; // 0x004a
	13'h0026: q3 = 16'h4c4d; // 0x004c
	13'h0027: q3 = 16'h4e4f; // 0x004e
	13'h0028: q3 = 16'h5051; // 0x0050
	13'h0029: q3 = 16'h5253; // 0x0052
	13'h002a: q3 = 16'h5455; // 0x0054
	13'h002b: q3 = 16'h5657; // 0x0056
	13'h002c: q3 = 16'h5859; // 0x0058
	13'h002d: q3 = 16'h5a5b; // 0x005a
	13'h002e: q3 = 16'h5c5d; // 0x005c
	13'h002f: q3 = 16'h5e5f; // 0x005e
	13'h0030: q3 = 16'h6061; // 0x0060
	13'h0031: q3 = 16'h6263; // 0x0062
	13'h0032: q3 = 16'h6465; // 0x0064
	13'h0033: q3 = 16'h6667; // 0x0066
	13'h0034: q3 = 16'h6869; // 0x0068
	13'h0035: q3 = 16'h6a6b; // 0x006a
	13'h0036: q3 = 16'h6c6d; // 0x006c
	13'h0037: q3 = 16'h6e6f; // 0x006e
	13'h0038: q3 = 16'h7071; // 0x0070
	13'h0039: q3 = 16'h7273; // 0x0072
	13'h003a: q3 = 16'h7475; // 0x0074
	13'h003b: q3 = 16'h7677; // 0x0076
	13'h003c: q3 = 16'h7879; // 0x0078
	13'h003d: q3 = 16'h7a7b; // 0x007a
	13'h003e: q3 = 16'h7c7d; // 0x007c
	13'h003f: q3 = 16'h7e7f; // 0x007e
	13'h0040: q3 = 16'h8081; // 0x0080
	13'h0041: q3 = 16'h8283; // 0x0082
	13'h0042: q3 = 16'h8485; // 0x0084
	13'h0043: q3 = 16'h8687; // 0x0086
	13'h0044: q3 = 16'h8889; // 0x0088
	13'h0045: q3 = 16'h8a8b; // 0x008a
	13'h0046: q3 = 16'h8c8d; // 0x008c
	13'h0047: q3 = 16'h8e8f; // 0x008e
	13'h0048: q3 = 16'h9091; // 0x0090
	13'h0049: q3 = 16'h9293; // 0x0092
	13'h004a: q3 = 16'h9495; // 0x0094
	13'h004b: q3 = 16'h9697; // 0x0096
	13'h004c: q3 = 16'h9899; // 0x0098
	13'h004d: q3 = 16'h9a9b; // 0x009a
	13'h004e: q3 = 16'h9c9d; // 0x009c
	13'h004f: q3 = 16'h9e9f; // 0x009e
	13'h0050: q3 = 16'ha0a1; // 0x00a0
	13'h0051: q3 = 16'ha2a3; // 0x00a2
	13'h0052: q3 = 16'ha4a5; // 0x00a4
	13'h0053: q3 = 16'ha6a7; // 0x00a6
	13'h0054: q3 = 16'ha8a9; // 0x00a8
	13'h0055: q3 = 16'haaab; // 0x00aa
	13'h0056: q3 = 16'hacad; // 0x00ac
	13'h0057: q3 = 16'haeaf; // 0x00ae
	13'h0058: q3 = 16'hb0b1; // 0x00b0
	13'h0059: q3 = 16'hb2b3; // 0x00b2
	13'h005a: q3 = 16'hb4b5; // 0x00b4
	13'h005b: q3 = 16'hb6b7; // 0x00b6
	13'h005c: q3 = 16'hb8b9; // 0x00b8
	13'h005d: q3 = 16'hbabb; // 0x00ba
	13'h005e: q3 = 16'hbcbd; // 0x00bc
	13'h005f: q3 = 16'hbebf; // 0x00be
	13'h0060: q3 = 16'hc0c1; // 0x00c0
	13'h0061: q3 = 16'hc2c3; // 0x00c2
	13'h0062: q3 = 16'hc4c5; // 0x00c4
	13'h0063: q3 = 16'hc6c7; // 0x00c6
	13'h0064: q3 = 16'hc8c9; // 0x00c8
	13'h0065: q3 = 16'hcacb; // 0x00ca
	13'h0066: q3 = 16'hcccd; // 0x00cc
	13'h0067: q3 = 16'hcecf; // 0x00ce
	13'h0068: q3 = 16'hd0d1; // 0x00d0
	13'h0069: q3 = 16'hd2d3; // 0x00d2
	13'h006a: q3 = 16'hd4d5; // 0x00d4
	13'h006b: q3 = 16'hd6d7; // 0x00d6
	13'h006c: q3 = 16'hd8d9; // 0x00d8
	13'h006d: q3 = 16'hdadb; // 0x00da
	13'h006e: q3 = 16'hdcdd; // 0x00dc
	13'h006f: q3 = 16'hdedf; // 0x00de
	13'h0070: q3 = 16'he0e1; // 0x00e0
	13'h0071: q3 = 16'he2e3; // 0x00e2
	13'h0072: q3 = 16'he4e5; // 0x00e4
	13'h0073: q3 = 16'he6e7; // 0x00e6
	13'h0074: q3 = 16'he8e9; // 0x00e8
	13'h0075: q3 = 16'heaeb; // 0x00ea
	13'h0076: q3 = 16'heced; // 0x00ec
	13'h0077: q3 = 16'heeef; // 0x00ee
	13'h0078: q3 = 16'hf0f1; // 0x00f0
	13'h0079: q3 = 16'hf2f3; // 0x00f2
	13'h007a: q3 = 16'hf4f5; // 0x00f4
	13'h007b: q3 = 16'hf6f7; // 0x00f6
	13'h007c: q3 = 16'hf8f9; // 0x00f8
	13'h007d: q3 = 16'hfafb; // 0x00fa
	13'h007e: q3 = 16'hfcfd; // 0x00fc
	13'h007f: q3 = 16'hfeff; // 0x00fe
	13'h0080: q3 = 16'h0000; // 0x0100
	13'h0081: q3 = 16'h000a; // 0x0102
	13'h0082: q3 = 16'h3000; // 0x0104
	13'h0083: q3 = 16'h011a; // 0x0106
	13'h0084: q3 = 16'h0117; // 0x0108
	13'h0085: q3 = 16'h000b; // 0x010a
	13'h0086: q3 = 16'h00a9; // 0x010c
	13'h0087: q3 = 16'h0085; // 0x010e
	13'h0088: q3 = 16'h002c; // 0x0110
	13'h0089: q3 = 16'h0060; // 0x0112
	13'h008a: q3 = 16'h004d; // 0x0114
	13'h008b: q3 = 16'h0021; // 0x0116
	13'h008c: q3 = 16'h0000; // 0x0118
	13'h008d: q3 = 16'h0000; // 0x011a
	13'h008e: q3 = 16'h0000; // 0x011c
	13'h008f: q3 = 16'h00c0; // 0x011e
	13'h0090: q3 = 16'h00c0; // 0x0120
	13'h0091: q3 = 16'h000a; // 0x0122
	13'h0092: q3 = 16'hffb8; // 0x0124
	13'h0093: q3 = 16'hffe8; // 0x0126
	13'h0094: q3 = 16'h004e; // 0x0128
	13'h0095: q3 = 16'h0000; // 0x012a
	13'h0096: q3 = 16'h011a; // 0x012c
	13'h0097: q3 = 16'h0000; // 0x012e
	13'h0098: q3 = 16'h0000; // 0x0130
	13'h0099: q3 = 16'h8136; // 0x0132
	13'h009a: q3 = 16'h0000; // 0x0134
	13'h009b: q3 = 16'hc106; // 0x0136
	13'h009c: q3 = 16'h0800; // 0x0138
	13'h009d: q3 = 16'h0000; // 0x013a
	13'h009e: q3 = 16'h0000; // 0x013c
	13'h009f: q3 = 16'h8136; // 0x013e
	13'h00a0: q3 = 16'h0000; // 0x0140
	13'h00a1: q3 = 16'hc11e; // 0x0142
	13'h00a2: q3 = 16'h0000; // 0x0144
	13'h00a3: q3 = 16'h0000; // 0x0146
	13'h00a4: q3 = 16'h0000; // 0x0148
	13'h00a5: q3 = 16'h0000; // 0x014a
	13'h00a6: q3 = 16'h00e0; // 0x014c
	13'h00a7: q3 = 16'h0000; // 0x014e
	13'h00a8: q3 = 16'h05d2; // 0x0150
	13'h00a9: q3 = 16'h0000; // 0x0152
	13'h00aa: q3 = 16'h0000; // 0x0154
	13'h00ab: q3 = 16'hc130; // 0x0156
	13'h00ac: q3 = 16'hffff; // 0x0158
	13'h00ad: q3 = 16'h0001; // 0x015a
	13'h00ae: q3 = 16'h0200; // 0x015c
	13'h00af: q3 = 16'h002a; // 0x015e
	13'h00b0: q3 = 16'haaaa; // 0x0160
	13'h00b1: q3 = 16'h0301; // 0x0162
	13'h00b2: q3 = 16'h0000; // 0x0164
	13'h00b3: q3 = 16'hc338; // 0x0166
	13'h00b4: q3 = 16'h0501; // 0x0168
	13'h00b5: q3 = 16'h0000; // 0x016a
	13'h00b6: q3 = 16'hc350; // 0x016c
	13'h00b7: q3 = 16'h8701; // 0x016e
	13'h00b8: q3 = 16'h0199; // 0x0170
	13'h00b9: q3 = 16'h0800; // 0x0172
	13'h00ba: q3 = 16'h8a01; // 0x0174
	13'h00bb: q3 = 16'h0800; // 0x0176
	13'h00bc: q3 = 16'h8701; // 0x0178
	13'h00bd: q3 = 16'h0199; // 0x017a
	13'h00be: q3 = 16'h0800; // 0x017c
	13'h00bf: q3 = 16'h8a01; // 0x017e
	13'h00c0: q3 = 16'h0800; // 0x0180
	13'h00c1: q3 = 16'h8701; // 0x0182
	13'h00c2: q3 = 16'h0199; // 0x0184
	13'h00c3: q3 = 16'h0800; // 0x0186
	13'h00c4: q3 = 16'h8a01; // 0x0188
	13'h00c5: q3 = 16'h1800; // 0x018a
	13'h00c6: q3 = 16'h0801; // 0x018c
	13'h00c7: q3 = 16'h0100; // 0x018e
	13'h00c8: q3 = 16'h0012; // 0x0190
	13'h00c9: q3 = 16'h1212; // 0x0192
	13'h00ca: q3 = 16'h1212; // 0x0194
	13'h00cb: q3 = 16'h1212; // 0x0196
	13'h00cc: q3 = 16'h1212; // 0x0198
	13'h00cd: q3 = 16'h1212; // 0x019a
	13'h00ce: q3 = 16'h1212; // 0x019c
	13'h00cf: q3 = 16'h1212; // 0x019e
	13'h00d0: q3 = 16'h0009; // 0x01a0
	13'h00d1: q3 = 16'h0d0e; // 0x01a2
	13'h00d2: q3 = 16'h0f10; // 0x01a4
	13'h00d3: q3 = 16'h1010; // 0x01a6
	13'h00d4: q3 = 16'h1111; // 0x01a8
	13'h00d5: q3 = 16'h1111; // 0x01aa
	13'h00d6: q3 = 16'h1111; // 0x01ac
	13'h00d7: q3 = 16'h1111; // 0x01ae
	13'h00d8: q3 = 16'h0005; // 0x01b0
	13'h00d9: q3 = 16'h090b; // 0x01b2
	13'h00da: q3 = 16'h0d0e; // 0x01b4
	13'h00db: q3 = 16'h0e0f; // 0x01b6
	13'h00dc: q3 = 16'h0f0f; // 0x01b8
	13'h00dd: q3 = 16'h1010; // 0x01ba
	13'h00de: q3 = 16'h1010; // 0x01bc
	13'h00df: q3 = 16'h1010; // 0x01be
	13'h00e0: q3 = 16'h0004; // 0x01c0
	13'h00e1: q3 = 16'h0709; // 0x01c2
	13'h00e2: q3 = 16'h0b0c; // 0x01c4
	13'h00e3: q3 = 16'h0d0d; // 0x01c6
	13'h00e4: q3 = 16'h0e0e; // 0x01c8
	13'h00e5: q3 = 16'h0f0f; // 0x01ca
	13'h00e6: q3 = 16'h0f0f; // 0x01cc
	13'h00e7: q3 = 16'h1010; // 0x01ce
	13'h00e8: q3 = 16'h0003; // 0x01d0
	13'h00e9: q3 = 16'h0507; // 0x01d2
	13'h00ea: q3 = 16'h090a; // 0x01d4
	13'h00eb: q3 = 16'h0b0c; // 0x01d6
	13'h00ec: q3 = 16'h0d0d; // 0x01d8
	13'h00ed: q3 = 16'h0e0e; // 0x01da
	13'h00ee: q3 = 16'h0e0f; // 0x01dc
	13'h00ef: q3 = 16'h0f0f; // 0x01de
	13'h00f0: q3 = 16'h0002; // 0x01e0
	13'h00f1: q3 = 16'h0406; // 0x01e2
	13'h00f2: q3 = 16'h0809; // 0x01e4
	13'h00f3: q3 = 16'h0a0b; // 0x01e6
	13'h00f4: q3 = 16'h0c0c; // 0x01e8
	13'h00f5: q3 = 16'h0d0d; // 0x01ea
	13'h00f6: q3 = 16'h0d0e; // 0x01ec
	13'h00f7: q3 = 16'h0e0e; // 0x01ee
	13'h00f8: q3 = 16'h0002; // 0x01f0
	13'h00f9: q3 = 16'h0405; // 0x01f2
	13'h00fa: q3 = 16'h0708; // 0x01f4
	13'h00fb: q3 = 16'h090a; // 0x01f6
	13'h00fc: q3 = 16'h0b0b; // 0x01f8
	13'h00fd: q3 = 16'h0c0c; // 0x01fa
	13'h00fe: q3 = 16'h0d0d; // 0x01fc
	13'h00ff: q3 = 16'h0d0e; // 0x01fe
	13'h0100: q3 = 16'h0002; // 0x0200
	13'h0101: q3 = 16'h0305; // 0x0202
	13'h0102: q3 = 16'h0607; // 0x0204
	13'h0103: q3 = 16'h0809; // 0x0206
	13'h0104: q3 = 16'h0a0a; // 0x0208
	13'h0105: q3 = 16'h0b0c; // 0x020a
	13'h0106: q3 = 16'h0c0c; // 0x020c
	13'h0107: q3 = 16'h0d0d; // 0x020e
	13'h0108: q3 = 16'h0001; // 0x0210
	13'h0109: q3 = 16'h0304; // 0x0212
	13'h010a: q3 = 16'h0506; // 0x0214
	13'h010b: q3 = 16'h0708; // 0x0216
	13'h010c: q3 = 16'h090a; // 0x0218
	13'h010d: q3 = 16'h0a0b; // 0x021a
	13'h010e: q3 = 16'h0b0c; // 0x021c
	13'h010f: q3 = 16'h0c0c; // 0x021e
	13'h0110: q3 = 16'h0001; // 0x0220
	13'h0111: q3 = 16'h0304; // 0x0222
	13'h0112: q3 = 16'h0506; // 0x0224
	13'h0113: q3 = 16'h0708; // 0x0226
	13'h0114: q3 = 16'h0809; // 0x0228
	13'h0115: q3 = 16'h0a0a; // 0x022a
	13'h0116: q3 = 16'h0b0b; // 0x022c
	13'h0117: q3 = 16'h0b0c; // 0x022e
	13'h0118: q3 = 16'h0001; // 0x0230
	13'h0119: q3 = 16'h0203; // 0x0232
	13'h011a: q3 = 16'h0405; // 0x0234
	13'h011b: q3 = 16'h0607; // 0x0236
	13'h011c: q3 = 16'h0808; // 0x0238
	13'h011d: q3 = 16'h090a; // 0x023a
	13'h011e: q3 = 16'h0a0a; // 0x023c
	13'h011f: q3 = 16'h0b0b; // 0x023e
	13'h0120: q3 = 16'h0001; // 0x0240
	13'h0121: q3 = 16'h0203; // 0x0242
	13'h0122: q3 = 16'h0405; // 0x0244
	13'h0123: q3 = 16'h0606; // 0x0246
	13'h0124: q3 = 16'h0708; // 0x0248
	13'h0125: q3 = 16'h0809; // 0x024a
	13'h0126: q3 = 16'h090a; // 0x024c
	13'h0127: q3 = 16'h0a0b; // 0x024e
	13'h0128: q3 = 16'h0001; // 0x0250
	13'h0129: q3 = 16'h0203; // 0x0252
	13'h012a: q3 = 16'h0405; // 0x0254
	13'h012b: q3 = 16'h0506; // 0x0256
	13'h012c: q3 = 16'h0707; // 0x0258
	13'h012d: q3 = 16'h0809; // 0x025a
	13'h012e: q3 = 16'h0909; // 0x025c
	13'h012f: q3 = 16'h0a0a; // 0x025e
	13'h0130: q3 = 16'h0001; // 0x0260
	13'h0131: q3 = 16'h0203; // 0x0262
	13'h0132: q3 = 16'h0304; // 0x0264
	13'h0133: q3 = 16'h0506; // 0x0266
	13'h0134: q3 = 16'h0607; // 0x0268
	13'h0135: q3 = 16'h0808; // 0x026a
	13'h0136: q3 = 16'h0909; // 0x026c
	13'h0137: q3 = 16'h090a; // 0x026e
	13'h0138: q3 = 16'h0001; // 0x0270
	13'h0139: q3 = 16'h0202; // 0x0272
	13'h013a: q3 = 16'h0304; // 0x0274
	13'h013b: q3 = 16'h0505; // 0x0276
	13'h013c: q3 = 16'h0607; // 0x0278
	13'h013d: q3 = 16'h0708; // 0x027a
	13'h013e: q3 = 16'h0809; // 0x027c
	13'h013f: q3 = 16'h0909; // 0x027e
	13'h0140: q3 = 16'h0001; // 0x0280
	13'h0141: q3 = 16'h0202; // 0x0282
	13'h0142: q3 = 16'h0304; // 0x0284
	13'h0143: q3 = 16'h0405; // 0x0286
	13'h0144: q3 = 16'h0606; // 0x0288
	13'h0145: q3 = 16'h0707; // 0x028a
	13'h0146: q3 = 16'h0808; // 0x028c
	13'h0147: q3 = 16'h0909; // 0x028e
	13'h0148: q3 = 16'hffcc; // 0x0290
	13'h0149: q3 = 16'hffda; // 0x0292
	13'h014a: q3 = 16'h0043; // 0x0294
	13'h014b: q3 = 16'hff82; // 0x0296
	13'h014c: q3 = 16'hffbd; // 0x0298
	13'h014d: q3 = 16'h0057; // 0x029a
	13'h014e: q3 = 16'hff5e; // 0x029c
	13'h014f: q3 = 16'hff7a; // 0x029e
	13'h0150: q3 = 16'h0026; // 0x02a0
	13'h0151: q3 = 16'h0000; // 0x02a2
	13'h0152: q3 = 16'h0000; // 0x02a4
	13'h0153: q3 = 16'h0000; // 0x02a6
	13'h0154: q3 = 16'h003c; // 0x02a8
	13'h0155: q3 = 16'h000c; // 0x02aa
	13'h0156: q3 = 16'h009c; // 0x02ac
	13'h0157: q3 = 16'hffa0; // 0x02ae
	13'h0158: q3 = 16'hffa0; // 0x02b0
	13'h0159: q3 = 16'h0014; // 0x02b2
	13'h015a: q3 = 16'h0000; // 0x02b4
	13'h015b: q3 = 16'hffcc; // 0x02b6
	13'h015c: q3 = 16'h0000; // 0x02b8
	13'h015d: q3 = 16'h0000; // 0x02ba
	13'h015e: q3 = 16'h8136; // 0x02bc
	13'h015f: q3 = 16'h0000; // 0x02be
	13'h0160: q3 = 16'hc290; // 0x02c0
	13'h0161: q3 = 16'h3500; // 0x02c2
	13'h0162: q3 = 16'h0000; // 0x02c4
	13'h0163: q3 = 16'h0000; // 0x02c6
	13'h0164: q3 = 16'h8136; // 0x02c8
	13'h0165: q3 = 16'h0000; // 0x02ca
	13'h0166: q3 = 16'hc2a8; // 0x02cc
	13'h0167: q3 = 16'h0000; // 0x02ce
	13'h0168: q3 = 16'h0000; // 0x02d0
	13'h0169: q3 = 16'h0000; // 0x02d2
	13'h016a: q3 = 16'h0000; // 0x02d4
	13'h016b: q3 = 16'h5859; // 0x02d6
	13'h016c: q3 = 16'h0000; // 0x02d8
	13'h016d: q3 = 16'h05dc; // 0x02da
	13'h016e: q3 = 16'h0000; // 0x02dc
	13'h016f: q3 = 16'h0000; // 0x02de
	13'h0170: q3 = 16'hc2ba; // 0x02e0
	13'h0171: q3 = 16'hffff; // 0x02e2
	13'h0172: q3 = 16'h0095; // 0x02e4
	13'h0173: q3 = 16'h8000; // 0x02e6
	13'h0174: q3 = 16'h000a; // 0x02e8
	13'h0175: q3 = 16'hbc25; // 0x02ea
	13'h0176: q3 = 16'h0000; // 0x02ec
	13'h0177: q3 = 16'h0030; // 0x02ee
	13'h0178: q3 = 16'h0080; // 0x02f0
	13'h0179: q3 = 16'h0080; // 0x02f2
	13'h017a: q3 = 16'h000a; // 0x02f4
	13'h017b: q3 = 16'hff90; // 0x02f6
	13'h017c: q3 = 16'hff90; // 0x02f8
	13'h017d: q3 = 16'h0008; // 0x02fa
	13'h017e: q3 = 16'h0000; // 0x02fc
	13'h017f: q3 = 16'h0000; // 0x02fe
	13'h0180: q3 = 16'h002d; // 0x0300
	13'h0181: q3 = 16'hffe4; // 0x0302
	13'h0182: q3 = 16'hfffa; // 0x0304
	13'h0183: q3 = 16'h0027; // 0x0306
	13'h0184: q3 = 16'hffec; // 0x0308
	13'h0185: q3 = 16'hffee; // 0x030a
	13'h0186: q3 = 16'h0007; // 0x030c
	13'h0187: q3 = 16'h0000; // 0x030e
	13'h0188: q3 = 16'h0000; // 0x0310
	13'h0189: q3 = 16'h7fff; // 0x0312
	13'h018a: q3 = 16'h0000; // 0x0314
	13'h018b: q3 = 16'h8136; // 0x0316
	13'h018c: q3 = 16'h0000; // 0x0318
	13'h018d: q3 = 16'hc2f0; // 0x031a
	13'h018e: q3 = 16'h0000; // 0x031c
	13'h018f: q3 = 16'h0000; // 0x031e
	13'h0190: q3 = 16'h0000; // 0x0320
	13'h0191: q3 = 16'h8136; // 0x0322
	13'h0192: q3 = 16'h0000; // 0x0324
	13'h0193: q3 = 16'hc30e; // 0x0326
	13'h0194: q3 = 16'h0000; // 0x0328
	13'h0195: q3 = 16'h0000; // 0x032a
	13'h0196: q3 = 16'hfff0; // 0x032c
	13'h0197: q3 = 16'hfff0; // 0x032e
	13'h0198: q3 = 16'h0020; // 0x0330
	13'h0199: q3 = 16'h0000; // 0x0332
	13'h019a: q3 = 16'h0000; // 0x0334
	13'h019b: q3 = 16'h7fff; // 0x0336
	13'h019c: q3 = 16'h0000; // 0x0338
	13'h019d: q3 = 16'h8136; // 0x033a
	13'h019e: q3 = 16'h0000; // 0x033c
	13'h019f: q3 = 16'hc32c; // 0x033e
	13'h01a0: q3 = 16'h0780; // 0x0340
	13'h01a1: q3 = 16'h0000; // 0x0342
	13'h01a2: q3 = 16'hffb6; // 0x0344
	13'h01a3: q3 = 16'hffd2; // 0x0346
	13'h01a4: q3 = 16'h001e; // 0x0348
	13'h01a5: q3 = 16'h0000; // 0x034a
	13'h01a6: q3 = 16'h0000; // 0x034c
	13'h01a7: q3 = 16'h7fff; // 0x034e
	13'h01a8: q3 = 16'h0000; // 0x0350
	13'h01a9: q3 = 16'h8136; // 0x0352
	13'h01aa: q3 = 16'h0000; // 0x0354
	13'h01ab: q3 = 16'hc344; // 0x0356
	13'h01ac: q3 = 16'h0580; // 0x0358
	13'h01ad: q3 = 16'h0000; // 0x035a
	13'h01ae: q3 = 16'h00b4; // 0x035c
	13'h01af: q3 = 16'h00ae; // 0x035e
	13'h01b0: q3 = 16'h000b; // 0x0360
	13'h01b1: q3 = 16'hffd0; // 0x0362
	13'h01b2: q3 = 16'hffd0; // 0x0364
	13'h01b3: q3 = 16'h0010; // 0x0366
	13'h01b4: q3 = 16'h0000; // 0x0368
	13'h01b5: q3 = 16'h0000; // 0x036a
	13'h01b6: q3 = 16'h7fff; // 0x036c
	13'h01b7: q3 = 16'h0000; // 0x036e
	13'h01b8: q3 = 16'h8136; // 0x0370
	13'h01b9: q3 = 16'h0000; // 0x0372
	13'h01ba: q3 = 16'hc35c; // 0x0374
	13'h01bb: q3 = 16'h0000; // 0x0376
	13'h01bc: q3 = 16'h0000; // 0x0378
	13'h01bd: q3 = 16'hffd0; // 0x037a
	13'h01be: q3 = 16'hffe8; // 0x037c
	13'h01bf: q3 = 16'h002f; // 0x037e
	13'h01c0: q3 = 16'h0000; // 0x0380
	13'h01c1: q3 = 16'h0000; // 0x0382
	13'h01c2: q3 = 16'h7fff; // 0x0384
	13'h01c3: q3 = 16'h0000; // 0x0386
	13'h01c4: q3 = 16'h8136; // 0x0388
	13'h01c5: q3 = 16'h0000; // 0x038a
	13'h01c6: q3 = 16'hc37a; // 0x038c
	13'h01c7: q3 = 16'h0480; // 0x038e
	13'h01c8: q3 = 16'h0000; // 0x0390
	13'h01c9: q3 = 16'h0001; // 0x0392
	13'h01ca: q3 = 16'h0200; // 0x0394
	13'h01cb: q3 = 16'h0038; // 0x0396
	13'h01cc: q3 = 16'he38e; // 0x0398
	13'h01cd: q3 = 16'h0301; // 0x039a
	13'h01ce: q3 = 16'h0000; // 0x039c
	13'h01cf: q3 = 16'hc338; // 0x039e
	13'h01d0: q3 = 16'h0501; // 0x03a0
	13'h01d1: q3 = 16'h0000; // 0x03a2
	13'h01d2: q3 = 16'hc350; // 0x03a4
	13'h01d3: q3 = 16'h8701; // 0x03a6
	13'h01d4: q3 = 16'h0445; // 0x03a8
	13'h01d5: q3 = 16'h03bb; // 0x03aa
	13'h01d6: q3 = 16'h8a01; // 0x03ac
	13'h01d7: q3 = 16'h019a; // 0x03ae
	13'h01d8: q3 = 16'h8701; // 0x03b0
	13'h01d9: q3 = 16'h0333; // 0x03b2
	13'h01da: q3 = 16'h03bc; // 0x03b4
	13'h01db: q3 = 16'h8a01; // 0x03b6
	13'h01dc: q3 = 16'h0199; // 0x03b8
	13'h01dd: q3 = 16'h8701; // 0x03ba
	13'h01de: q3 = 16'h028a; // 0x03bc
	13'h01df: q3 = 16'h03bc; // 0x03be
	13'h01e0: q3 = 16'h8a01; // 0x03c0
	13'h01e1: q3 = 16'h019a; // 0x03c2
	13'h01e2: q3 = 16'h8701; // 0x03c4
	13'h01e3: q3 = 16'h0222; // 0x03c6
	13'h01e4: q3 = 16'h0777; // 0x03c8
	13'h01e5: q3 = 16'h8a01; // 0x03ca
	13'h01e6: q3 = 16'h0333; // 0x03cc
	13'h01e7: q3 = 16'h8701; // 0x03ce
	13'h01e8: q3 = 16'h028a; // 0x03d0
	13'h01e9: q3 = 16'h03bc; // 0x03d2
	13'h01ea: q3 = 16'h8a01; // 0x03d4
	13'h01eb: q3 = 16'h019a; // 0x03d6
	13'h01ec: q3 = 16'h8701; // 0x03d8
	13'h01ed: q3 = 16'h0222; // 0x03da
	13'h01ee: q3 = 16'h1666; // 0x03dc
	13'h01ef: q3 = 16'h8a01; // 0x03de
	13'h01f0: q3 = 16'h099a; // 0x03e0
	13'h01f1: q3 = 16'h0801; // 0x03e2
	13'h01f2: q3 = 16'h0100; // 0x03e4
	13'h01f3: q3 = 16'hff80; // 0x03e6
	13'h01f4: q3 = 16'hff80; // 0x03e8
	13'h01f5: q3 = 16'h0010; // 0x03ea
	13'h01f6: q3 = 16'h0110; // 0x03ec
	13'h01f7: q3 = 16'h0108; // 0x03ee
	13'h01f8: q3 = 16'h001f; // 0x03f0
	13'h01f9: q3 = 16'h0000; // 0x03f2
	13'h01fa: q3 = 16'h0000; // 0x03f4
	13'h01fb: q3 = 16'h0000; // 0x03f6
	13'h01fc: q3 = 16'h0040; // 0x03f8
	13'h01fd: q3 = 16'h0040; // 0x03fa
	13'h01fe: q3 = 16'h0010; // 0x03fc
	13'h01ff: q3 = 16'hffd4; // 0x03fe
	13'h0200: q3 = 16'hffdd; // 0x0400
	13'h0201: q3 = 16'h001d; // 0x0402
	13'h0202: q3 = 16'h0000; // 0x0404
	13'h0203: q3 = 16'hff80; // 0x0406
	13'h0204: q3 = 16'h0000; // 0x0408
	13'h0205: q3 = 16'h0080; // 0x040a
	13'h0206: q3 = 16'h0038; // 0x040c
	13'h0207: q3 = 16'h00e0; // 0x040e
	13'h0208: q3 = 16'h0000; // 0x0410
	13'h0209: q3 = 16'h0000; // 0x0412
	13'h020a: q3 = 16'h8136; // 0x0414
	13'h020b: q3 = 16'h0000; // 0x0416
	13'h020c: q3 = 16'hc3e6; // 0x0418
	13'h020d: q3 = 16'h0800; // 0x041a
	13'h020e: q3 = 16'h0000; // 0x041c
	13'h020f: q3 = 16'h0000; // 0x041e
	13'h0210: q3 = 16'h8136; // 0x0420
	13'h0211: q3 = 16'h0000; // 0x0422
	13'h0212: q3 = 16'hc3f8; // 0x0424
	13'h0213: q3 = 16'h0000; // 0x0426
	13'h0214: q3 = 16'h0000; // 0x0428
	13'h0215: q3 = 16'h0000; // 0x042a
	13'h0216: q3 = 16'hc40a; // 0x042c
	13'h0217: q3 = 16'h00e0; // 0x042e
	13'h0218: q3 = 16'h0000; // 0x0430
	13'h0219: q3 = 16'h0000; // 0x0432
	13'h021a: q3 = 16'h0000; // 0x0434
	13'h021b: q3 = 16'h0009; // 0x0436
	13'h021c: q3 = 16'h0063; // 0x0438
	13'h021d: q3 = 16'h0055; // 0x043a
	13'h021e: q3 = 16'h002a; // 0x043c
	13'h021f: q3 = 16'h0000; // 0x043e
	13'h0220: q3 = 16'h0014; // 0x0440
	13'h0221: q3 = 16'h0000; // 0x0442
	13'h0222: q3 = 16'h0061; // 0x0444
	13'h0223: q3 = 16'h005b; // 0x0446
	13'h0224: q3 = 16'h000e; // 0x0448
	13'h0225: q3 = 16'hffce; // 0x044a
	13'h0226: q3 = 16'hffd7; // 0x044c
	13'h0227: q3 = 16'h001f; // 0x044e
	13'h0228: q3 = 16'h0000; // 0x0450
	13'h0229: q3 = 16'h0080; // 0x0452
	13'h022a: q3 = 16'h0000; // 0x0454
	13'h022b: q3 = 16'h0000; // 0x0456
	13'h022c: q3 = 16'h8136; // 0x0458
	13'h022d: q3 = 16'h0000; // 0x045a
	13'h022e: q3 = 16'hc432; // 0x045c
	13'h022f: q3 = 16'h0800; // 0x045e
	13'h0230: q3 = 16'h0000; // 0x0460
	13'h0231: q3 = 16'h0000; // 0x0462
	13'h0232: q3 = 16'h8136; // 0x0464
	13'h0233: q3 = 16'h0000; // 0x0466
	13'h0234: q3 = 16'hc444; // 0x0468
	13'h0235: q3 = 16'h0000; // 0x046a
	13'h0236: q3 = 16'h0000; // 0x046c
	13'h0237: q3 = 16'h0000; // 0x046e
	13'h0238: q3 = 16'h0000; // 0x0470
	13'h0239: q3 = 16'h6c6d; // 0x0472
	13'h023a: q3 = 16'h0000; // 0x0474
	13'h023b: q3 = 16'h0040; // 0x0476
	13'h023c: q3 = 16'h00c2; // 0x0478
	13'h023d: q3 = 16'h0000; // 0x047a
	13'h023e: q3 = 16'h0000; // 0x047c
	13'h023f: q3 = 16'h0000; // 0x047e
	13'h0240: q3 = 16'hc476; // 0x0480
	13'h0241: q3 = 16'h0000; // 0x0482
	13'h0242: q3 = 16'h0000; // 0x0484
	13'h0243: q3 = 16'h03e8; // 0x0486
	13'h0244: q3 = 16'h0001; // 0x0488
	13'h0245: q3 = 16'h0000; // 0x048a
	13'h0246: q3 = 16'hc412; // 0x048c
	13'h0247: q3 = 16'h0000; // 0x048e
	13'h0248: q3 = 16'hc47e; // 0x0490
	13'h0249: q3 = 16'h0000; // 0x0492
	13'h024a: q3 = 16'h0000; // 0x0494
	13'h024b: q3 = 16'hc456; // 0x0496
	13'h024c: q3 = 16'hffff; // 0x0498
	13'h024d: q3 = 16'h0000; // 0x049a
	13'h024e: q3 = 16'h0000; // 0x049c
	13'h024f: q3 = 16'h0000; // 0x049e
	13'h0250: q3 = 16'hffa7; // 0x04a0
	13'h0251: q3 = 16'hffab; // 0x04a2
	13'h0252: q3 = 16'h000c; // 0x04a4
	13'h0253: q3 = 16'hffda; // 0x04a6
	13'h0254: q3 = 16'hfff3; // 0x04a8
	13'h0255: q3 = 16'h0043; // 0x04aa
	13'h0256: q3 = 16'h0000; // 0x04ac
	13'h0257: q3 = 16'h0000; // 0x04ae
	13'h0258: q3 = 16'h0000; // 0x04b0
	13'h0259: q3 = 16'h00c0; // 0x04b2
	13'h025a: q3 = 16'h005a; // 0x04b4
	13'h025b: q3 = 16'h00e0; // 0x04b6
	13'h025c: q3 = 16'h0000; // 0x04b8
	13'h025d: q3 = 16'h0000; // 0x04ba
	13'h025e: q3 = 16'h8136; // 0x04bc
	13'h025f: q3 = 16'h0000; // 0x04be
	13'h0260: q3 = 16'hc49a; // 0x04c0
	13'h0261: q3 = 16'h0e00; // 0x04c2
	13'h0262: q3 = 16'h0000; // 0x04c4
	13'h0263: q3 = 16'h0000; // 0x04c6
	13'h0264: q3 = 16'h8136; // 0x04c8
	13'h0265: q3 = 16'h0000; // 0x04ca
	13'h0266: q3 = 16'hc4a0; // 0x04cc
	13'h0267: q3 = 16'h0780; // 0x04ce
	13'h0268: q3 = 16'h0000; // 0x04d0
	13'h0269: q3 = 16'h0000; // 0x04d2
	13'h026a: q3 = 16'hc4b2; // 0x04d4
	13'h026b: q3 = 16'h00e0; // 0x04d6
	13'h026c: q3 = 16'h0000; // 0x04d8
	13'h026d: q3 = 16'h0000; // 0x04da
	13'h026e: q3 = 16'h0000; // 0x04dc
	13'h026f: q3 = 16'h0000; // 0x04de
	13'h0270: q3 = 16'hffb5; // 0x04e0
	13'h0271: q3 = 16'hffb7; // 0x04e2
	13'h0272: q3 = 16'h000e; // 0x04e4
	13'h0273: q3 = 16'hffc0; // 0x04e6
	13'h0274: q3 = 16'hfff3; // 0x04e8
	13'h0275: q3 = 16'h0041; // 0x04ea
	13'h0276: q3 = 16'h0000; // 0x04ec
	13'h0277: q3 = 16'h00c0; // 0x04ee
	13'h0278: q3 = 16'h0000; // 0x04f0
	13'h0279: q3 = 16'h0060; // 0x04f2
	13'h027a: q3 = 16'h0060; // 0x04f4
	13'h027b: q3 = 16'h00e0; // 0x04f6
	13'h027c: q3 = 16'h0000; // 0x04f8
	13'h027d: q3 = 16'h0000; // 0x04fa
	13'h027e: q3 = 16'h8136; // 0x04fc
	13'h027f: q3 = 16'h0000; // 0x04fe
	13'h0280: q3 = 16'hc4da; // 0x0500
	13'h0281: q3 = 16'h0000; // 0x0502
	13'h0282: q3 = 16'h0000; // 0x0504
	13'h0283: q3 = 16'h0000; // 0x0506
	13'h0284: q3 = 16'h8136; // 0x0508
	13'h0285: q3 = 16'h0000; // 0x050a
	13'h0286: q3 = 16'hc4e0; // 0x050c
	13'h0287: q3 = 16'h0780; // 0x050e
	13'h0288: q3 = 16'h0000; // 0x0510
	13'h0289: q3 = 16'h0000; // 0x0512
	13'h028a: q3 = 16'hc4f2; // 0x0514
	13'h028b: q3 = 16'h00e0; // 0x0516
	13'h028c: q3 = 16'h0000; // 0x0518
	13'h028d: q3 = 16'h0040; // 0x051a
	13'h028e: q3 = 16'h0059; // 0x051c
	13'h028f: q3 = 16'h0000; // 0x051e
	13'h0290: q3 = 16'h0000; // 0x0520
	13'h0291: q3 = 16'h0000; // 0x0522
	13'h0292: q3 = 16'hc51a; // 0x0524
	13'h0293: q3 = 16'h0000; // 0x0526
	13'h0294: q3 = 16'h0000; // 0x0528
	13'h0295: q3 = 16'h0040; // 0x052a
	13'h0296: q3 = 16'h0057; // 0x052c
	13'h0297: q3 = 16'h0000; // 0x052e
	13'h0298: q3 = 16'h0000; // 0x0530
	13'h0299: q3 = 16'h0000; // 0x0532
	13'h029a: q3 = 16'hc52a; // 0x0534
	13'h029b: q3 = 16'h0000; // 0x0536
	13'h029c: q3 = 16'h0000; // 0x0538
	13'h029d: q3 = 16'h0fa0; // 0x053a
	13'h029e: q3 = 16'h0001; // 0x053c
	13'h029f: q3 = 16'h0000; // 0x053e
	13'h02a0: q3 = 16'hc4ba; // 0x0540
	13'h02a1: q3 = 16'h0000; // 0x0542
	13'h02a2: q3 = 16'hc522; // 0x0544
	13'h02a3: q3 = 16'h0001; // 0x0546
	13'h02a4: q3 = 16'h0000; // 0x0548
	13'h02a5: q3 = 16'hc4fa; // 0x054a
	13'h02a6: q3 = 16'h0000; // 0x054c
	13'h02a7: q3 = 16'hc4fa; // 0x054e
	13'h02a8: q3 = 16'hffff; // 0x0550
	13'h02a9: q3 = 16'h0094; // 0x0552
	13'h02aa: q3 = 16'h8000; // 0x0554
	13'h02ab: q3 = 16'h2020; // 0x0556
	13'h02ac: q3 = 16'h2020; // 0x0558
	13'h02ad: q3 = 16'h11f6; // 0x055a
	13'h02ae: q3 = 16'hf50f; // 0x055c
	13'h02af: q3 = 16'h2020; // 0x055e
	13'h02b0: q3 = 16'hf712; // 0x0560
	13'h02b1: q3 = 16'hf1f1; // 0x0562
	13'h02b2: q3 = 16'hf1f1; // 0x0564
	13'h02b3: q3 = 16'h2015; // 0x0566
	13'h02b4: q3 = 16'h13f1; // 0x0568
	13'h02b5: q3 = 16'hf1f1; // 0x056a
	13'h02b6: q3 = 16'hf1f1; // 0x056c
	13'h02b7: q3 = 16'h2014; // 0x056e
	13'h02b8: q3 = 16'hf1f1; // 0x0570
	13'h02b9: q3 = 16'hf1f1; // 0x0572
	13'h02ba: q3 = 16'hf1f1; // 0x0574
	13'h02bb: q3 = 16'h2016; // 0x0576
	13'h02bc: q3 = 16'hf1f1; // 0x0578
	13'h02bd: q3 = 16'hf1f1; // 0x057a
	13'h02be: q3 = 16'hf1f1; // 0x057c
	13'h02bf: q3 = 16'h2017; // 0x057e
	13'h02c0: q3 = 16'hf1f1; // 0x0580
	13'h02c1: q3 = 16'hf1f1; // 0x0582
	13'h02c2: q3 = 16'hf1f1; // 0x0584
	13'h02c3: q3 = 16'h20f8; // 0x0586
	13'h02c4: q3 = 16'h18f1; // 0x0588
	13'h02c5: q3 = 16'hf1f1; // 0x058a
	13'h02c6: q3 = 16'hf1f1; // 0x058c
	13'h02c7: q3 = 16'h2020; // 0x058e
	13'h02c8: q3 = 16'hf9fd; // 0x0590
	13'h02c9: q3 = 16'hf1f1; // 0x0592
	13'h02ca: q3 = 16'hf1f1; // 0x0594
	13'h02cb: q3 = 16'h2020; // 0x0596
	13'h02cc: q3 = 16'h2020; // 0x0598
	13'h02cd: q3 = 16'hfaff; // 0x059a
	13'h02ce: q3 = 16'h10fc; // 0x059c
	13'h02cf: q3 = 16'h2020; // 0x059e
	13'h02d0: q3 = 16'h2020; // 0x05a0
	13'h02d1: q3 = 16'h7ef5; // 0x05a2
	13'h02d2: q3 = 16'h607c; // 0x05a4
	13'h02d3: q3 = 16'h2020; // 0x05a6
	13'h02d4: q3 = 16'hf712; // 0x05a8
	13'h02d5: q3 = 16'hf1f1; // 0x05aa
	13'h02d6: q3 = 16'hf175; // 0x05ac
	13'h02d7: q3 = 16'h2020; // 0x05ae
	13'h02d8: q3 = 16'h13f1; // 0x05b0
	13'h02d9: q3 = 16'hf1f1; // 0x05b2
	13'h02da: q3 = 16'hf176; // 0x05b4
	13'h02db: q3 = 16'h2014; // 0x05b6
	13'h02dc: q3 = 16'hf1f1; // 0x05b8
	13'h02dd: q3 = 16'hf1f1; // 0x05ba
	13'h02de: q3 = 16'hf177; // 0x05bc
	13'h02df: q3 = 16'h2016; // 0x05be
	13'h02e0: q3 = 16'hf1f1; // 0x05c0
	13'h02e1: q3 = 16'hf1f1; // 0x05c2
	13'h02e2: q3 = 16'hf178; // 0x05c4
	13'h02e3: q3 = 16'h2017; // 0x05c6
	13'h02e4: q3 = 16'hf1f1; // 0x05c8
	13'h02e5: q3 = 16'hf1f1; // 0x05ca
	13'h02e6: q3 = 16'hf179; // 0x05cc
	13'h02e7: q3 = 16'h2020; // 0x05ce
	13'h02e8: q3 = 16'h18f1; // 0x05d0
	13'h02e9: q3 = 16'hf1f1; // 0x05d2
	13'h02ea: q3 = 16'hf17a; // 0x05d4
	13'h02eb: q3 = 16'h2020; // 0x05d6
	13'h02ec: q3 = 16'hfbfd; // 0x05d8
	13'h02ed: q3 = 16'hf1f1; // 0x05da
	13'h02ee: q3 = 16'hf17b; // 0x05dc
	13'h02ef: q3 = 16'h2020; // 0x05de
	13'h02f0: q3 = 16'h2020; // 0x05e0
	13'h02f1: q3 = 16'h7f10; // 0x05e2
	13'h02f2: q3 = 16'h617d; // 0x05e4
	13'h02f3: q3 = 16'h2020; // 0x05e6
	13'h02f4: q3 = 16'h207e; // 0x05e8
	13'h02f5: q3 = 16'hf50f; // 0x05ea
	13'h02f6: q3 = 16'h8963; // 0x05ec
	13'h02f7: q3 = 16'h20f7; // 0x05ee
	13'h02f8: q3 = 16'h12f1; // 0x05f0
	13'h02f9: q3 = 16'hf1f1; // 0x05f2
	13'h02fa: q3 = 16'h7580; // 0x05f4
	13'h02fb: q3 = 16'h1513; // 0x05f6
	13'h02fc: q3 = 16'hf1f1; // 0x05f8
	13'h02fd: q3 = 16'hf1f1; // 0x05fa
	13'h02fe: q3 = 16'h7681; // 0x05fc
	13'h02ff: q3 = 16'h14f1; // 0x05fe
	13'h0300: q3 = 16'hf1f1; // 0x0600
	13'h0301: q3 = 16'hf1f1; // 0x0602
	13'h0302: q3 = 16'h7782; // 0x0604
	13'h0303: q3 = 16'h16f1; // 0x0606
	13'h0304: q3 = 16'hf1f1; // 0x0608
	13'h0305: q3 = 16'hf1f1; // 0x060a
	13'h0306: q3 = 16'h7883; // 0x060c
	13'h0307: q3 = 16'h17f1; // 0x060e
	13'h0308: q3 = 16'hf1f1; // 0x0610
	13'h0309: q3 = 16'hf1f1; // 0x0612
	13'h030a: q3 = 16'h7984; // 0x0614
	13'h030b: q3 = 16'hfe18; // 0x0616
	13'h030c: q3 = 16'hf1f1; // 0x0618
	13'h030d: q3 = 16'hf1f1; // 0x061a
	13'h030e: q3 = 16'h7a85; // 0x061c
	13'h030f: q3 = 16'h20f9; // 0x061e
	13'h0310: q3 = 16'hfdf1; // 0x0620
	13'h0311: q3 = 16'hf1f1; // 0x0622
	13'h0312: q3 = 16'h7b86; // 0x0624
	13'h0313: q3 = 16'h2020; // 0x0626
	13'h0314: q3 = 16'h207f; // 0x0628
	13'h0315: q3 = 16'h10fc; // 0x062a
	13'h0316: q3 = 16'h8887; // 0x062c
	13'h0317: q3 = 16'h66bf; // 0x062e
	13'h0318: q3 = 16'h15a7; // 0x0630
	13'h0319: q3 = 16'hb92f; // 0x0632
	13'h031a: q3 = 16'h3b8e; // 0x0634
	13'h031b: q3 = 16'h3e47; // 0x0636
	13'h031c: q3 = 16'h14ad; // 0x0638
	13'h031d: q3 = 16'h0254; // 0x063a
	13'h031e: q3 = 16'h5914; // 0x063c
	13'h031f: q3 = 16'h2143; // 0x063e
	13'h0320: q3 = 16'h1b44; // 0x0640
	13'h0321: q3 = 16'h0a51; // 0x0642
	13'h0322: q3 = 16'h0141; // 0x0644
	13'h0323: q3 = 16'h5002; // 0x0646
	13'h0324: q3 = 16'h1141; // 0x0648
	13'h0325: q3 = 16'h0941; // 0x064a
	13'h0326: q3 = 16'h0000; // 0x064c
	13'h0327: q3 = 16'h157c; // 0x064e
	13'h0328: q3 = 16'h0000; // 0x0650
	13'h0329: q3 = 16'h1588; // 0x0652
	13'h032a: q3 = 16'h0000; // 0x0654
	13'h032b: q3 = 16'h1592; // 0x0656
	13'h032c: q3 = 16'h0000; // 0x0658
	13'h032d: q3 = 16'h15a2; // 0x065a
	13'h032e: q3 = 16'h0000; // 0x065c
	13'h032f: q3 = 16'h15b2; // 0x065e
	13'h0330: q3 = 16'h0000; // 0x0660
	13'h0331: q3 = 16'h15ba; // 0x0662
	13'h0332: q3 = 16'h0000; // 0x0664
	13'h0333: q3 = 16'h15c2; // 0x0666
	13'h0334: q3 = 16'h0000; // 0x0668
	13'h0335: q3 = 16'h15ca; // 0x066a
	13'h0336: q3 = 16'h0000; // 0x066c
	13'h0337: q3 = 16'h15d2; // 0x066e
	13'h0338: q3 = 16'h0000; // 0x0670
	13'h0339: q3 = 16'h15da; // 0x0672
	13'h033a: q3 = 16'h0003; // 0x0674
	13'h033b: q3 = 16'h0200; // 0x0676
	13'h033c: q3 = 16'h004f; // 0x0678
	13'h033d: q3 = 16'ha4fa; // 0x067a
	13'h033e: q3 = 16'h0303; // 0x067c
	13'h033f: q3 = 16'h0000; // 0x067e
	13'h0340: q3 = 16'hf332; // 0x0680
	13'h0341: q3 = 16'h0000; // 0x0682
	13'h0342: q3 = 16'hc36e; // 0x0684
	13'h0343: q3 = 16'h0503; // 0x0686
	13'h0344: q3 = 16'h0000; // 0x0688
	13'h0345: q3 = 16'hf34a; // 0x068a
	13'h0346: q3 = 16'h0000; // 0x068c
	13'h0347: q3 = 16'hc386; // 0x068e
	13'h0348: q3 = 16'h8703; // 0x0690
	13'h0349: q3 = 16'h0333; // 0x0692
	13'h034a: q3 = 16'h0666; // 0x0694
	13'h034b: q3 = 16'h0800; // 0x0696
	13'h034c: q3 = 16'h0701; // 0x0698
	13'h034d: q3 = 16'h0222; // 0x069a
	13'h034e: q3 = 16'h8a02; // 0x069c
	13'h034f: q3 = 16'h0800; // 0x069e
	13'h0350: q3 = 16'h8703; // 0x06a0
	13'h0351: q3 = 16'h0199; // 0x06a2
	13'h0352: q3 = 16'h0445; // 0x06a4
	13'h0353: q3 = 16'h0800; // 0x06a6
	13'h0354: q3 = 16'h0701; // 0x06a8
	13'h0355: q3 = 16'h01b1; // 0x06aa
	13'h0356: q3 = 16'h8a02; // 0x06ac
	13'h0357: q3 = 16'h0800; // 0x06ae
	13'h0358: q3 = 16'h8702; // 0x06b0
	13'h0359: q3 = 16'h05b3; // 0x06b2
	13'h035a: q3 = 16'h0800; // 0x06b4
	13'h035b: q3 = 16'h0701; // 0x06b6
	13'h035c: q3 = 16'h0222; // 0x06b8
	13'h035d: q3 = 16'h8a02; // 0x06ba
	13'h035e: q3 = 16'h0800; // 0x06bc
	13'h035f: q3 = 16'h8703; // 0x06be
	13'h0360: q3 = 16'h01b1; // 0x06c0
	13'h0361: q3 = 16'h0445; // 0x06c2
	13'h0362: q3 = 16'h0800; // 0x06c4
	13'h0363: q3 = 16'h0701; // 0x06c6
	13'h0364: q3 = 16'h016c; // 0x06c8
	13'h0365: q3 = 16'h8a02; // 0x06ca
	13'h0366: q3 = 16'h0800; // 0x06cc
	13'h0367: q3 = 16'h8703; // 0x06ce
	13'h0368: q3 = 16'h0199; // 0x06d0
	13'h0369: q3 = 16'h0333; // 0x06d2
	13'h036a: q3 = 16'h0800; // 0x06d4
	13'h036b: q3 = 16'h8a02; // 0x06d6
	13'h036c: q3 = 16'h0800; // 0x06d8
	13'h036d: q3 = 16'h8702; // 0x06da
	13'h036e: q3 = 16'h0445; // 0x06dc
	13'h036f: q3 = 16'h0800; // 0x06de
	13'h0370: q3 = 16'h8a02; // 0x06e0
	13'h0371: q3 = 16'h0800; // 0x06e2
	13'h0372: q3 = 16'h8702; // 0x06e4
	13'h0373: q3 = 16'h0333; // 0x06e6
	13'h0374: q3 = 16'h0800; // 0x06e8
	13'h0375: q3 = 16'h8a03; // 0x06ea
	13'h0376: q3 = 16'h0800; // 0x06ec
	13'h0377: q3 = 16'h0803; // 0x06ee
	13'h0378: q3 = 16'h0100; // 0x06f0
	13'h0379: q3 = 16'h0005; // 0x06f2
	13'h037a: q3 = 16'h0200; // 0x06f4
	13'h037b: q3 = 16'h0033; // 0x06f6
	13'h037c: q3 = 16'h3333; // 0x06f8
	13'h037d: q3 = 16'h0305; // 0x06fa
	13'h037e: q3 = 16'h0000; // 0x06fc
	13'h037f: q3 = 16'hf332; // 0x06fe
	13'h0380: q3 = 16'h0000; // 0x0700
	13'h0381: q3 = 16'hc314; // 0x0702
	13'h0382: q3 = 16'h0505; // 0x0704
	13'h0383: q3 = 16'h0000; // 0x0706
	13'h0384: q3 = 16'hf34a; // 0x0708
	13'h0385: q3 = 16'h0000; // 0x070a
	13'h0386: q3 = 16'hc320; // 0x070c
	13'h0387: q3 = 16'h8705; // 0x070e
	13'h0388: q3 = 16'h0199; // 0x0710
	13'h0389: q3 = 16'h0666; // 0x0712
	13'h038a: q3 = 16'h0400; // 0x0714
	13'h038b: q3 = 16'h8a05; // 0x0716
	13'h038c: q3 = 16'h0400; // 0x0718
	13'h038d: q3 = 16'h8705; // 0x071a
	13'h038e: q3 = 16'h01e7; // 0x071c
	13'h038f: q3 = 16'h088b; // 0x071e
	13'h0390: q3 = 16'h0400; // 0x0720
	13'h0391: q3 = 16'h8a05; // 0x0722
	13'h0392: q3 = 16'h0400; // 0x0724
	13'h0393: q3 = 16'h8705; // 0x0726
	13'h0394: q3 = 16'h0222; // 0x0728
	13'h0395: q3 = 16'h079c; // 0x072a
	13'h0396: q3 = 16'h0400; // 0x072c
	13'h0397: q3 = 16'h0701; // 0x072e
	13'h0398: q3 = 16'h01e7; // 0x0730
	13'h0399: q3 = 16'h8a04; // 0x0732
	13'h039a: q3 = 16'h0400; // 0x0734
	13'h039b: q3 = 16'h0704; // 0x0736
	13'h039c: q3 = 16'h06c7; // 0x0738
	13'h039d: q3 = 16'h8a01; // 0x073a
	13'h039e: q3 = 16'h0400; // 0x073c
	13'h039f: q3 = 16'h0701; // 0x073e
	13'h03a0: q3 = 16'h0199; // 0x0740
	13'h03a1: q3 = 16'h8a04; // 0x0742
	13'h03a2: q3 = 16'h0400; // 0x0744
	13'h03a3: q3 = 16'h8704; // 0x0746
	13'h03a4: q3 = 16'h0666; // 0x0748
	13'h03a5: q3 = 16'h0400; // 0x074a
	13'h03a6: q3 = 16'h8a04; // 0x074c
	13'h03a7: q3 = 16'h0400; // 0x074e
	13'h03a8: q3 = 16'h0601; // 0x0750
	13'h03a9: q3 = 16'h0479; // 0x0752
	13'h03aa: q3 = 16'hfb9a; // 0x0754
	13'h03ab: q3 = 16'h8b01; // 0x0756
	13'h03ac: q3 = 16'h0333; // 0x0758
	13'h03ad: q3 = 16'h0800; // 0x075a
	13'h03ae: q3 = 16'h8704; // 0x075c
	13'h03af: q3 = 16'h0ccc; // 0x075e
	13'h03b0: q3 = 16'h0400; // 0x0760
	13'h03b1: q3 = 16'h8a04; // 0x0762
	13'h03b2: q3 = 16'h0400; // 0x0764
	13'h03b3: q3 = 16'h8a01; // 0x0766
	13'h03b4: q3 = 16'h0800; // 0x0768
	13'h03b5: q3 = 16'h8804; // 0x076a
	13'h03b6: q3 = 16'h1000; // 0x076c
	13'h03b7: q3 = 16'h0801; // 0x076e
	13'h03b8: q3 = 16'h0100; // 0x0770
	13'h03b9: q3 = 16'h00ac; // 0x0772
	13'h03ba: q3 = 16'h00aa; // 0x0774
	13'h03bb: q3 = 16'h0003; // 0x0776
	13'h03bc: q3 = 16'hff00; // 0x0778
	13'h03bd: q3 = 16'hff00; // 0x077a
	13'h03be: q3 = 16'h0006; // 0x077c
	13'h03bf: q3 = 16'hfed0; // 0x077e
	13'h03c0: q3 = 16'hfed8; // 0x0780
	13'h03c1: q3 = 16'h0013; // 0x0782
	13'h03c2: q3 = 16'h0000; // 0x0784
	13'h03c3: q3 = 16'h0000; // 0x0786
	13'h03c4: q3 = 16'h0000; // 0x0788
	13'h03c5: q3 = 16'h0078; // 0x078a
	13'h03c6: q3 = 16'h0071; // 0x078c
	13'h03c7: q3 = 16'h0009; // 0x078e
	13'h03c8: q3 = 16'hffa0; // 0x0790
	13'h03c9: q3 = 16'hffa0; // 0x0792
	13'h03ca: q3 = 16'h0014; // 0x0794
	13'h03cb: q3 = 16'h0000; // 0x0796
	13'h03cc: q3 = 16'h00ac; // 0x0798
	13'h03cd: q3 = 16'h0000; // 0x079a
	13'h03ce: q3 = 16'h0000; // 0x079c
	13'h03cf: q3 = 16'h8136; // 0x079e
	13'h03d0: q3 = 16'h0000; // 0x07a0
	13'h03d1: q3 = 16'hc772; // 0x07a2
	13'h03d2: q3 = 16'h1c00; // 0x07a4
	13'h03d3: q3 = 16'h0000; // 0x07a6
	13'h03d4: q3 = 16'h0000; // 0x07a8
	13'h03d5: q3 = 16'h8136; // 0x07aa
	13'h03d6: q3 = 16'h0000; // 0x07ac
	13'h03d7: q3 = 16'hc78a; // 0x07ae
	13'h03d8: q3 = 16'h0380; // 0x07b0
	13'h03d9: q3 = 16'h0000; // 0x07b2
	13'h03da: q3 = 16'h0000; // 0x07b4
	13'h03db: q3 = 16'h0000; // 0x07b6
	13'h03dc: q3 = 16'h00e0; // 0x07b8
	13'h03dd: q3 = 16'h0000; // 0x07ba
	13'h03de: q3 = 16'h0640; // 0x07bc
	13'h03df: q3 = 16'h0000; // 0x07be
	13'h03e0: q3 = 16'h0000; // 0x07c0
	13'h03e1: q3 = 16'hc79c; // 0x07c2
	13'h03e2: q3 = 16'hffff; // 0x07c4
	13'h03e3: q3 = 16'h001a; // 0x07c6
	13'h03e4: q3 = 16'h0004; // 0x07c8
	13'h03e5: q3 = 16'h000e; // 0x07ca
	13'h03e6: q3 = 16'h000a; // 0x07cc
	13'h03e7: q3 = 16'h0004; // 0x07ce
	13'h03e8: q3 = 16'h0095; // 0x07d0
	13'h03e9: q3 = 16'h4000; // 0x07d2
	13'h03ea: q3 = 16'h0090; // 0x07d4
	13'h03eb: q3 = 16'h0000; // 0x07d6
	13'h03ec: q3 = 16'h0004; // 0x07d8
	13'h03ed: q3 = 16'h0000; // 0x07da
	13'h03ee: q3 = 16'h0095; // 0x07dc
	13'h03ef: q3 = 16'h8000; // 0x07de
	13'h03f0: q3 = 16'h0094; // 0x07e0
	13'h03f1: q3 = 16'h8000; // 0x07e2
	13'h03f2: q3 = 16'h0090; // 0x07e4
	13'h03f3: q3 = 16'h0000; // 0x07e6
	13'h03f4: q3 = 16'h0000; // 0x07e8
	13'h03f5: q3 = 16'hc150; // 0x07ea
	13'h03f6: q3 = 16'h0000; // 0x07ec
	13'h03f7: q3 = 16'hf56e; // 0x07ee
	13'h03f8: q3 = 16'h0000; // 0x07f0
	13'h03f9: q3 = 16'he05e; // 0x07f2
	13'h03fa: q3 = 16'h0000; // 0x07f4
	13'h03fb: q3 = 16'hfed4; // 0x07f6
	13'h03fc: q3 = 16'h0006; // 0x07f8
	13'h03fd: q3 = 16'h000c; // 0x07fa
	13'h03fe: q3 = 16'h0004; // 0x07fc
	13'h03ff: q3 = 16'h0002; // 0x07fe
	13'h0400: q3 = 16'h0003; // 0x0800
	13'h0401: q3 = 16'h0019; // 0x0802
	13'h0402: q3 = 16'h0012; // 0x0804
	13'h0403: q3 = 16'h000b; // 0x0806
	13'h0404: q3 = 16'h000e; // 0x0808
	13'h0405: q3 = 16'h0014; // 0x080a
	13'h0406: q3 = 16'h0001; // 0x080c
	13'h0407: q3 = 16'h05b6; // 0x080e
	13'h0408: q3 = 16'h0000; // 0x0810
	13'h0409: q3 = 16'h2718; // 0x0812
	13'h040a: q3 = 16'h0000; // 0x0814
	13'h040b: q3 = 16'h2728; // 0x0816
	13'h040c: q3 = 16'h0000; // 0x0818
	13'h040d: q3 = 16'h2736; // 0x081a
	13'h040e: q3 = 16'h0000; // 0x081c
	13'h040f: q3 = 16'h274e; // 0x081e
	13'h0410: q3 = 16'h0000; // 0x0820
	13'h0411: q3 = 16'h275e; // 0x0822
	13'h0412: q3 = 16'h0000; // 0x0824
	13'h0413: q3 = 16'h27aa; // 0x0826
	13'h0414: q3 = 16'h0000; // 0x0828
	13'h0415: q3 = 16'h27c8; // 0x082a
	13'h0416: q3 = 16'h0000; // 0x082c
	13'h0417: q3 = 16'h27e2; // 0x082e
	13'h0418: q3 = 16'h0000; // 0x0830
	13'h0419: q3 = 16'hc2da; // 0x0832
	13'h041a: q3 = 16'h0000; // 0x0834
	13'h041b: q3 = 16'hf5c2; // 0x0836
	13'h041c: q3 = 16'h0000; // 0x0838
	13'h041d: q3 = 16'he0d6; // 0x083a
	13'h041e: q3 = 16'h0000; // 0x083c
	13'h041f: q3 = 16'hff22; // 0x083e
	13'h0420: q3 = 16'h0000; // 0x0840
	13'h0421: q3 = 16'h2b58; // 0x0842
	13'h0422: q3 = 16'h0000; // 0x0844
	13'h0423: q3 = 16'h2b5e; // 0x0846
	13'h0424: q3 = 16'h0000; // 0x0848
	13'h0425: q3 = 16'h2b80; // 0x084a
	13'h0426: q3 = 16'h0000; // 0x084c
	13'h0427: q3 = 16'h2b92; // 0x084e
	13'h0428: q3 = 16'h0004; // 0x0850
	13'h0429: q3 = 16'h0078; // 0x0852
	13'h042a: q3 = 16'h0005; // 0x0854
	13'h042b: q3 = 16'h0001; // 0x0856
	13'h042c: q3 = 16'h0090; // 0x0858
	13'h042d: q3 = 16'h0003; // 0x085a
	13'h042e: q3 = 16'h0002; // 0x085c
	13'h042f: q3 = 16'h0060; // 0x085e
	13'h0430: q3 = 16'h0006; // 0x0860
	13'h0431: q3 = 16'h0003; // 0x0862
	13'h0432: q3 = 16'h0080; // 0x0864
	13'h0433: q3 = 16'h0004; // 0x0866
	13'h0434: q3 = 16'h0002; // 0x0868
	13'h0435: q3 = 16'h0060; // 0x086a
	13'h0436: q3 = 16'h0006; // 0x086c
	13'h0437: q3 = 16'h0001; // 0x086e
	13'h0438: q3 = 16'h0090; // 0x0870
	13'h0439: q3 = 16'h0003; // 0x0872
	13'h043a: q3 = 16'h0003; // 0x0874
	13'h043b: q3 = 16'h0080; // 0x0876
	13'h043c: q3 = 16'h0004; // 0x0878
	13'h043d: q3 = 16'h0004; // 0x087a
	13'h043e: q3 = 16'h0078; // 0x087c
	13'h043f: q3 = 16'h0005; // 0x087e
	13'h0440: q3 = 16'hc0c1; // 0x0880
	13'h0441: q3 = 16'hc2c1; // 0x0882
	13'h0442: q3 = 16'h672d; // 0x0884
	13'h0443: q3 = 16'h2e30; // 0x0886
	13'h0444: q3 = 16'h3030; // 0x0888
	13'h0445: q3 = 16'h3030; // 0x088a
	13'h0446: q3 = 16'h3030; // 0x088c
	13'h0447: q3 = 16'h3000; // 0x088e
	13'h0448: q3 = 16'h6060; // 0x0890
	13'h0449: q3 = 16'h602f; // 0x0892
	13'h044a: q3 = 16'h3630; // 0x0894
	13'h044b: q3 = 16'h3030; // 0x0896
	13'h044c: q3 = 16'h3030; // 0x0898
	13'h044d: q3 = 16'h3000; // 0x089a
	13'h044e: q3 = 16'h6f6f; // 0x089c
	13'h044f: q3 = 16'h6f6f; // 0x089e
	13'h0450: q3 = 16'h6f6f; // 0x08a0
	13'h0451: q3 = 16'h191a; // 0x08a2
	13'h0452: q3 = 16'h3030; // 0x08a4
	13'h0453: q3 = 16'h3070; // 0x08a6
	13'h0454: q3 = 16'h7070; // 0x08a8
	13'h0455: q3 = 16'h7070; // 0x08aa
	13'h0456: q3 = 16'h7038; // 0x08ac
	13'h0457: q3 = 16'h393a; // 0x08ae
	13'h0458: q3 = 16'h3b30; // 0x08b0
	13'h0459: q3 = 16'h7171; // 0x08b2
	13'h045a: q3 = 16'h7171; // 0x08b4
	13'h045b: q3 = 16'h7171; // 0x08b6
	13'h045c: q3 = 16'h3c3d; // 0x08b8
	13'h045d: q3 = 16'h3e3f; // 0x08ba
	13'h045e: q3 = 16'h3072; // 0x08bc
	13'h045f: q3 = 16'h7272; // 0x08be
	13'h0460: q3 = 16'h7272; // 0x08c0
	13'h0461: q3 = 16'h721b; // 0x08c2
	13'h0462: q3 = 16'h3730; // 0x08c4
	13'h0463: q3 = 16'h3030; // 0x08c6
	13'h0464: q3 = 16'h0016; // 0x08c8
	13'h0465: q3 = 16'h0011; // 0x08ca
	13'h0466: q3 = 16'h000d; // 0x08cc
	13'h0467: q3 = 16'h000a; // 0x08ce
	13'h0468: q3 = 16'h0008; // 0x08d0
	13'h0469: q3 = 16'h0000; // 0x08d2
	13'h046a: q3 = 16'h0000; // 0x08d4
	13'h046b: q3 = 16'h0000; // 0x08d6
	13'h046c: q3 = 16'h0000; // 0x08d8
	13'h046d: q3 = 16'h0101; // 0x08da
	13'h046e: q3 = 16'h0514; // 0x08dc
	13'h046f: q3 = 16'h0101; // 0x08de
	13'h0470: q3 = 16'h0100; // 0x08e0
	13'h0471: q3 = 16'h0000; // 0x08e2
	13'h0472: q3 = 16'h0010; // 0x08e4
	13'h0473: q3 = 16'h0010; // 0x08e6
	13'h0474: q3 = 16'h0060; // 0x08e8
	13'h0475: q3 = 16'h0042; // 0x08ea
	13'h0476: q3 = 16'h002b; // 0x08ec
	13'h0477: q3 = 16'h003b; // 0x08ee
	13'h0478: q3 = 16'h0112; // 0x08f0
	13'h0479: q3 = 16'h010e; // 0x08f2
	13'h047a: q3 = 16'h0012; // 0x08f4
	13'h047b: q3 = 16'h5300; // 0x08f6
	13'h047c: q3 = 16'h5300; // 0x08f8
	13'h047d: q3 = 16'h0001; // 0x08fa
	13'h047e: q3 = 16'h0000; // 0x08fc
	13'h047f: q3 = 16'h0000; // 0x08fe
	13'h0480: q3 = 16'h0000; // 0x0900
	13'h0481: q3 = 16'h0076; // 0x0902
	13'h0482: q3 = 16'h006a; // 0x0904
	13'h0483: q3 = 16'h0012; // 0x0906
	13'h0484: q3 = 16'hff98; // 0x0908
	13'h0485: q3 = 16'hfff6; // 0x090a
	13'h0486: q3 = 16'h009d; // 0x090c
	13'h0487: q3 = 16'hff00; // 0x090e
	13'h0488: q3 = 16'hff00; // 0x0910
	13'h0489: q3 = 16'h0001; // 0x0912
	13'h048a: q3 = 16'h0500; // 0x0914
	13'h048b: q3 = 16'h0500; // 0x0916
	13'h048c: q3 = 16'h0001; // 0x0918
	13'h048d: q3 = 16'hffd0; // 0x091a
	13'h048e: q3 = 16'hffd6; // 0x091c
	13'h048f: q3 = 16'h0009; // 0x091e
	13'h0490: q3 = 16'hffdf; // 0x0920
	13'h0491: q3 = 16'hfff7; // 0x0922
	13'h0492: q3 = 16'h0028; // 0x0924
	13'h0493: q3 = 16'hffd4; // 0x0926
	13'h0494: q3 = 16'hffe6; // 0x0928
	13'h0495: q3 = 16'h0013; // 0x092a
	13'h0496: q3 = 16'h0000; // 0x092c
	13'h0497: q3 = 16'h0010; // 0x092e
	13'h0498: q3 = 16'h0000; // 0x0930
	13'h0499: q3 = 16'h00e0; // 0x0932
	13'h049a: q3 = 16'h00b0; // 0x0934
	13'h049b: q3 = 16'h0000; // 0x0936
	13'h049c: q3 = 16'h004f; // 0x0938
	13'h049d: q3 = 16'h00e0; // 0x093a
	13'h049e: q3 = 16'h0000; // 0x093c
	13'h049f: q3 = 16'h0000; // 0x093e
	13'h04a0: q3 = 16'h8136; // 0x0940
	13'h04a1: q3 = 16'h0000; // 0x0942
	13'h04a2: q3 = 16'hc8e4; // 0x0944
	13'h04a3: q3 = 16'h0900; // 0x0946
	13'h04a4: q3 = 16'h0000; // 0x0948
	13'h04a5: q3 = 16'h0000; // 0x094a
	13'h04a6: q3 = 16'h8136; // 0x094c
	13'h04a7: q3 = 16'h0000; // 0x094e
	13'h04a8: q3 = 16'hc902; // 0x0950
	13'h04a9: q3 = 16'h0000; // 0x0952
	13'h04aa: q3 = 16'h0000; // 0x0954
	13'h04ab: q3 = 16'h0000; // 0x0956
	13'h04ac: q3 = 16'hc932; // 0x0958
	13'h04ad: q3 = 16'h00e0; // 0x095a
	13'h04ae: q3 = 16'h0000; // 0x095c
	13'h04af: q3 = 16'h0000; // 0x095e
	13'h04b0: q3 = 16'h00b0; // 0x0960
	13'h04b1: q3 = 16'h0040; // 0x0962
	13'h04b2: q3 = 16'h004f; // 0x0964
	13'h04b3: q3 = 16'h0000; // 0x0966
	13'h04b4: q3 = 16'h0000; // 0x0968
	13'h04b5: q3 = 16'h0000; // 0x096a
	13'h04b6: q3 = 16'hc95e; // 0x096c
	13'h04b7: q3 = 16'h0000; // 0x096e
	13'h04b8: q3 = 16'h0000; // 0x0970
	13'h04b9: q3 = 16'h07d0; // 0x0972
	13'h04ba: q3 = 16'h0001; // 0x0974
	13'h04bb: q3 = 16'h0000; // 0x0976
	13'h04bc: q3 = 16'hc93e; // 0x0978
	13'h04bd: q3 = 16'h0000; // 0x097a
	13'h04be: q3 = 16'hc96a; // 0x097c
	13'h04bf: q3 = 16'hffff; // 0x097e
	13'h04c0: q3 = 16'h0080; // 0x0980
	13'h04c1: q3 = 16'h0000; // 0x0982
	13'h04c2: q3 = 16'h0080; // 0x0984
	13'h04c3: q3 = 16'h0000; // 0x0986
	13'h04c4: q3 = 16'h0004; // 0x0988
	13'h04c5: q3 = 16'h0005; // 0x098a
	13'h04c6: q3 = 16'h0006; // 0x098c
	13'h04c7: q3 = 16'h0007; // 0x098e
	13'h04c8: q3 = 16'h0400; // 0x0990
	13'h04c9: q3 = 16'h0500; // 0x0992
	13'h04ca: q3 = 16'h0600; // 0x0994
	13'h04cb: q3 = 16'h0700; // 0x0996
	13'h04cc: q3 = 16'h0089; // 0x0998
	13'h04cd: q3 = 16'h0086; // 0x099a
	13'h04ce: q3 = 16'h00c9; // 0x099c
	13'h04cf: q3 = 16'h00c6; // 0x099e
	13'h04d0: q3 = 16'h0000; // 0x09a0
	13'h04d1: q3 = 16'h00c4; // 0x09a2
	13'h04d2: q3 = 16'h0000; // 0x09a4
	13'h04d3: q3 = 16'h00c5; // 0x09a6
	13'h04d4: q3 = 16'h0000; // 0x09a8
	13'h04d5: q3 = 16'h00c4; // 0x09aa
	13'h04d6: q3 = 16'h0000; // 0x09ac
	13'h04d7: q3 = 16'h00c5; // 0x09ae
	13'h04d8: q3 = 16'h0000; // 0x09b0
	13'h04d9: q3 = 16'h0000; // 0x09b2
	13'h04da: q3 = 16'h0040; // 0x09b4
	13'h04db: q3 = 16'h0040; // 0x09b6
	13'h04dc: q3 = 16'h00c0; // 0x09b8
	13'h04dd: q3 = 16'h0080; // 0x09ba
	13'h04de: q3 = 16'h0080; // 0x09bc
	13'h04df: q3 = 16'h0000; // 0x09be
	13'h04e0: q3 = 16'h0013; // 0x09c0
	13'h04e1: q3 = 16'h001a; // 0x09c2
	13'h04e2: q3 = 16'h001b; // 0x09c4
	13'h04e3: q3 = 16'h0001; // 0x09c6
	13'h04e4: q3 = 16'h001c; // 0x09c8
	13'h04e5: q3 = 16'h0000; // 0x09ca
	13'h04e6: q3 = 16'h0016; // 0x09cc
	13'h04e7: q3 = 16'h0180; // 0x09ce
	13'h04e8: q3 = 16'h0030; // 0x09d0
	13'h04e9: q3 = 16'h0001; // 0x09d2
	13'h04ea: q3 = 16'h000a; // 0x09d4
	13'h04eb: q3 = 16'h0200; // 0x09d6
	13'h04ec: q3 = 16'h0020; // 0x09d8
	13'h04ed: q3 = 16'h0004; // 0x09da
	13'h04ee: q3 = 16'h0011; // 0x09dc
	13'h04ef: q3 = 16'h0240; // 0x09de
	13'h04f0: q3 = 16'h0010; // 0x09e0
	13'h04f1: q3 = 16'h0002; // 0x09e2
	13'h04f2: q3 = 16'h000f; // 0x09e4
	13'h04f3: q3 = 16'h0240; // 0x09e6
	13'h04f4: q3 = 16'h0040; // 0x09e8
	13'h04f5: q3 = 16'h0035; // 0x09ea
	13'h04f6: q3 = 16'h0018; // 0x09ec
	13'h04f7: q3 = 16'h0180; // 0x09ee
	13'h04f8: q3 = 16'h00ff; // 0x09f0
	13'h04f9: q3 = 16'h040f; // 0x09f2
	13'h04fa: q3 = 16'h1621; // 0x09f4
	13'h04fb: q3 = 16'h2833; // 0x09f6
	13'h04fc: q3 = 16'h3a45; // 0x09f8
	13'h04fd: q3 = 16'h4800; // 0x09fa
	13'h04fe: q3 = 16'hcf85; // 0x09fc
	13'h04ff: q3 = 16'h0185; // 0x09fe
	13'h0500: q3 = 16'hcf85; // 0x0a00
	13'h0501: q3 = 16'h0185; // 0x0a02
	13'h0502: q3 = 16'h0000; // 0x0a04
	13'h0503: q3 = 16'h0080; // 0x0a06
	13'h0504: q3 = 16'h80c0; // 0x0a08
	13'h0505: q3 = 16'h4040; // 0x0a0a
	13'h0506: q3 = 16'h3030; // 0x0a0c
	13'h0507: q3 = 16'h0000; // 0x0a0e
	13'h0508: q3 = 16'h2056; // 0x0a10
	13'h0509: q3 = 16'h4f52; // 0x0a12
	13'h050a: q3 = 16'h4245; // 0x0a14
	13'h050b: q3 = 16'h4900; // 0x0a16
	13'h050c: q3 = 16'h0606; // 0x0a18
	13'h050d: q3 = 16'h0505; // 0x0a1a
	13'h050e: q3 = 16'h0504; // 0x0a1c
	13'h050f: q3 = 16'h0404; // 0x0a1e
	13'h0510: q3 = 16'h0303; // 0x0a20
	13'h0511: q3 = 16'h0302; // 0x0a22
	13'h0512: q3 = 16'h0202; // 0x0a24
	13'h0513: q3 = 16'h0101; // 0x0a26
	13'h0514: q3 = 16'h0100; // 0x0a28
	13'h0515: q3 = 16'h0000; // 0x0a2a
	13'h0516: q3 = 16'h0101; // 0x0a2c
	13'h0517: q3 = 16'h0102; // 0x0a2e
	13'h0518: q3 = 16'h0202; // 0x0a30
	13'h0519: q3 = 16'h0303; // 0x0a32
	13'h051a: q3 = 16'h0304; // 0x0a34
	13'h051b: q3 = 16'h0404; // 0x0a36
	13'h051c: q3 = 16'h0505; // 0x0a38
	13'h051d: q3 = 16'h0506; // 0x0a3a
	13'h051e: q3 = 16'h0606; // 0x0a3c
	13'h051f: q3 = 16'h0707; // 0x0a3e
	13'h0520: q3 = 16'h0708; // 0x0a40
	13'h0521: q3 = 16'h0808; // 0x0a42
	13'h0522: q3 = 16'h0909; // 0x0a44
	13'h0523: q3 = 16'h090a; // 0x0a46
	13'h0524: q3 = 16'h0a0a; // 0x0a48
	13'h0525: q3 = 16'h0b0b; // 0x0a4a
	13'h0526: q3 = 16'h0b0c; // 0x0a4c
	13'h0527: q3 = 16'h0c0c; // 0x0a4e
	13'h0528: q3 = 16'h0b0b; // 0x0a50
	13'h0529: q3 = 16'h0b0a; // 0x0a52
	13'h052a: q3 = 16'h0a0a; // 0x0a54
	13'h052b: q3 = 16'h0909; // 0x0a56
	13'h052c: q3 = 16'h0908; // 0x0a58
	13'h052d: q3 = 16'h0808; // 0x0a5a
	13'h052e: q3 = 16'h0707; // 0x0a5c
	13'h052f: q3 = 16'h0706; // 0x0a5e
	13'h0530: q3 = 16'h0000; // 0x0a60
	13'h0531: q3 = 16'h0020; // 0x0a62
	13'h0532: q3 = 16'h0040; // 0x0a64
	13'h0533: q3 = 16'h0060; // 0x0a66
	13'h0534: q3 = 16'hffff; // 0x0a68
	13'h0535: q3 = 16'h00a8; // 0x0a6a
	13'h0536: q3 = 16'h00c8; // 0x0a6c
	13'h0537: q3 = 16'h00e8; // 0x0a6e
	13'h0538: q3 = 16'h0108; // 0x0a70
	13'h0539: q3 = 16'hffff; // 0x0a72
	13'h053a: q3 = 16'h0150; // 0x0a74
	13'h053b: q3 = 16'h0170; // 0x0a76
	13'h053c: q3 = 16'h0190; // 0x0a78
	13'h053d: q3 = 16'h01b0; // 0x0a7a
	13'h053e: q3 = 16'hffff; // 0x0a7c
	13'h053f: q3 = 16'h0080; // 0x0a7e
	13'h0540: q3 = 16'h0088; // 0x0a80
	13'h0541: q3 = 16'h0090; // 0x0a82
	13'h0542: q3 = 16'h0098; // 0x0a84
	13'h0543: q3 = 16'h00a0; // 0x0a86
	13'h0544: q3 = 16'h0128; // 0x0a88
	13'h0545: q3 = 16'h0130; // 0x0a8a
	13'h0546: q3 = 16'h0138; // 0x0a8c
	13'h0547: q3 = 16'h0140; // 0x0a8e
	13'h0548: q3 = 16'h0148; // 0x0a90
	13'h0549: q3 = 16'h01d0; // 0x0a92
	13'h054a: q3 = 16'h01d8; // 0x0a94
	13'h054b: q3 = 16'h01e0; // 0x0a96
	13'h054c: q3 = 16'h01e8; // 0x0a98
	13'h054d: q3 = 16'h01f0; // 0x0a9a
	13'h054e: q3 = 16'h00d8; // 0x0a9c
	13'h054f: q3 = 16'h0105; // 0x0a9e
	13'h0550: q3 = 16'h0106; // 0x0aa0
	13'h0551: q3 = 16'h0107; // 0x0aa2
	13'h0552: q3 = 16'h0108; // 0x0aa4
	13'h0553: q3 = 16'h0109; // 0x0aa6
	13'h0554: q3 = 16'h010a; // 0x0aa8
	13'h0555: q3 = 16'h010b; // 0x0aaa
	13'h0556: q3 = 16'h010c; // 0x0aac
	13'h0557: q3 = 16'h010d; // 0x0aae
	13'h0558: q3 = 16'h010e; // 0x0ab0
	13'h0559: q3 = 16'h000f; // 0x0ab2
	13'h055a: q3 = 16'h0006; // 0x0ab4
	13'h055b: q3 = 16'h0003; // 0x0ab6
	13'h055c: q3 = 16'h0003; // 0x0ab8
	13'h055d: q3 = 16'h0002; // 0x0aba
	13'h055e: q3 = 16'h0002; // 0x0abc
	13'h055f: q3 = 16'h0002; // 0x0abe
	13'h0560: q3 = 16'h0001; // 0x0ac0
	13'h0561: q3 = 16'h0001; // 0x0ac2
	13'h0562: q3 = 16'h0002; // 0x0ac4
	13'h0563: q3 = 16'h0004; // 0x0ac6
	13'h0564: q3 = 16'h00e9; // 0x0ac8
	13'h0565: q3 = 16'h00ea; // 0x0aca
	13'h0566: q3 = 16'h00eb; // 0x0acc
	13'h0567: q3 = 16'h0100; // 0x0ace
	13'h0568: q3 = 16'h0101; // 0x0ad0
	13'h0569: q3 = 16'h0102; // 0x0ad2
	13'h056a: q3 = 16'h0103; // 0x0ad4
	13'h056b: q3 = 16'h0104; // 0x0ad6
	13'h056c: q3 = 16'h0040; // 0x0ad8
	13'h056d: q3 = 16'h00e1; // 0x0ada
	13'h056e: q3 = 16'h00e2; // 0x0adc
	13'h056f: q3 = 16'h00e3; // 0x0ade
	13'h0570: q3 = 16'h00e4; // 0x0ae0
	13'h0571: q3 = 16'h00e5; // 0x0ae2
	13'h0572: q3 = 16'h00e6; // 0x0ae4
	13'h0573: q3 = 16'h00e7; // 0x0ae6
	13'h0574: q3 = 16'h00e8; // 0x0ae8
	13'h0575: q3 = 16'h0040; // 0x0aea
	13'h0576: q3 = 16'h00d9; // 0x0aec
	13'h0577: q3 = 16'h00da; // 0x0aee
	13'h0578: q3 = 16'h00db; // 0x0af0
	13'h0579: q3 = 16'h00dc; // 0x0af2
	13'h057a: q3 = 16'h00dd; // 0x0af4
	13'h057b: q3 = 16'h00de; // 0x0af6
	13'h057c: q3 = 16'h00df; // 0x0af8
	13'h057d: q3 = 16'h00e0; // 0x0afa
	13'h057e: q3 = 16'h0040; // 0x0afc
	13'h057f: q3 = 16'h0002; // 0x0afe
	13'h0580: q3 = 16'heb2c; // 0x0b00
	13'h0581: q3 = 16'h0001; // 0x0b02
	13'h0582: q3 = 16'h07ac; // 0x0b04
	13'h0583: q3 = 16'h0000; // 0x0b06
	13'h0584: q3 = 16'h0000; // 0x0b08
	13'h0585: q3 = 16'h0013; // 0x0b0a
	13'h0586: q3 = 16'h001a; // 0x0b0c
	13'h0587: q3 = 16'h001b; // 0x0b0e
	13'h0588: q3 = 16'h0001; // 0x0b10
	13'h0589: q3 = 16'h001c; // 0x0b12
	13'h058a: q3 = 16'h0000; // 0x0b14
	13'h058b: q3 = 16'h0000; // 0x0b16
	13'h058c: q3 = 16'h0054; // 0x0b18
	13'h058d: q3 = 16'hd72c; // 0x0b1a
	13'h058e: q3 = 16'h002b; // 0x0b1c
	13'h058f: q3 = 16'h2f8a; // 0x0b1e
	13'h0590: q3 = 16'h2000; // 0x0b20
	13'h0591: q3 = 16'hbf09; // 0x0b22
	13'h0592: q3 = 16'h0a0b; // 0x0b24
	13'h0593: q3 = 16'h2030; // 0x0b26
	13'h0594: q3 = 16'h3030; // 0x0b28
	13'h0595: q3 = 16'h3030; // 0x0b2a
	13'h0596: q3 = 16'h3000; // 0x0b2c
	13'h0597: q3 = 16'h8c8c; // 0x0b2e
	13'h0598: q3 = 16'h8c8c; // 0x0b30
	13'h0599: q3 = 16'h8c8c; // 0x0b32
	13'h059a: q3 = 16'h2122; // 0x0b34
	13'h059b: q3 = 16'h2324; // 0x0b36
	13'h059c: q3 = 16'h3000; // 0x0b38
	13'h059d: q3 = 16'hcccc; // 0x0b3a
	13'h059e: q3 = 16'hcccc; // 0x0b3c
	13'h059f: q3 = 16'hcccc; // 0x0b3e
	13'h05a0: q3 = 16'h8182; // 0x0b40
	13'h05a1: q3 = 16'h8384; // 0x0b42
	13'h05a2: q3 = 16'h3000; // 0x0b44
	13'h05a3: q3 = 16'hbe1c; // 0x0b46
	13'h05a4: q3 = 16'h1d1e; // 0x0b48
	13'h05a5: q3 = 16'h1f30; // 0x0b4a
	13'h05a6: q3 = 16'h3030; // 0x0b4c
	13'h05a7: q3 = 16'h3030; // 0x0b4e
	13'h05a8: q3 = 16'h3000; // 0x0b50
	13'h05a9: q3 = 16'hfafb; // 0x0b52
	13'h05aa: q3 = 16'hfcfd; // 0x0b54
	13'h05ab: q3 = 16'hfeba; // 0x0b56
	13'h05ac: q3 = 16'hbbbb; // 0x0b58
	13'h05ad: q3 = 16'h2526; // 0x0b5a
	13'h05ae: q3 = 16'h2728; // 0x0b5c
	13'h05af: q3 = 16'h292a; // 0x0b5e
	13'h05b0: q3 = 16'h2bf9; // 0x0b60
	13'h05b1: q3 = 16'h7374; // 0x0b62
	13'h05b2: q3 = 16'h7576; // 0x0b64
	13'h05b3: q3 = 16'h7778; // 0x0b66
	13'h05b4: q3 = 16'h797a; // 0x0b68
	13'h05b5: q3 = 16'h7b7c; // 0x0b6a
	13'h05b6: q3 = 16'h7d7e; // 0x0b6c
	13'h05b7: q3 = 16'h8000; // 0x0b6e
	13'h05b8: q3 = 16'h3030; // 0x0b70
	13'h05b9: q3 = 16'h0000; // 0x0b72
	13'h05ba: q3 = 16'h4041; // 0x0b74
	13'h05bb: q3 = 16'h42c7; // 0x0b76
	13'h05bc: q3 = 16'hcacd; // 0x0b78
	13'h05bd: q3 = 16'hd0d3; // 0x0b7a
	13'h05be: q3 = 16'hd6d9; // 0x0b7c
	13'h05bf: q3 = 16'hd9d9; // 0x0b7e
	13'h05c0: q3 = 16'hd9d9; // 0x0b80
	13'h05c1: q3 = 16'hd6d3; // 0x0b82
	13'h05c2: q3 = 16'hd0cd; // 0x0b84
	13'h05c3: q3 = 16'hcac7; // 0x0b86
	13'h05c4: q3 = 16'h4241; // 0x0b88
	13'h05c5: q3 = 16'h4000; // 0x0b8a
	13'h05c6: q3 = 16'h3030; // 0x0b8c
	13'h05c7: q3 = 16'h3030; // 0x0b8e
	13'h05c8: q3 = 16'h3030; // 0x0b90
	13'h05c9: q3 = 16'h8f92; // 0x0b92
	13'h05ca: q3 = 16'h9598; // 0x0b94
	13'h05cb: q3 = 16'h9b9e; // 0x0b96
	13'h05cc: q3 = 16'ha1a4; // 0x0b98
	13'h05cd: q3 = 16'ha7aa; // 0x0b9a
	13'h05ce: q3 = 16'hadb0; // 0x0b9c
	13'h05cf: q3 = 16'hb330; // 0x0b9e
	13'h05d0: q3 = 16'h3030; // 0x0ba0
	13'h05d1: q3 = 16'h3000; // 0x0ba2
	13'h05d2: q3 = 16'h5151; // 0x0ba4
	13'h05d3: q3 = 16'h5252; // 0x0ba6
	13'h05d4: q3 = 16'h5253; // 0x0ba8
	13'h05d5: q3 = 16'h5455; // 0x0baa
	13'h05d6: q3 = 16'h5657; // 0x0bac
	13'h05d7: q3 = 16'h5757; // 0x0bae
	13'h05d8: q3 = 16'h5757; // 0x0bb0
	13'h05d9: q3 = 16'h5655; // 0x0bb2
	13'h05da: q3 = 16'h5453; // 0x0bb4
	13'h05db: q3 = 16'h5252; // 0x0bb6
	13'h05dc: q3 = 16'h5251; // 0x0bb8
	13'h05dd: q3 = 16'h5100; // 0x0bba
	13'h05de: q3 = 16'h0001; // 0x0bbc
	13'h05df: q3 = 16'h0008; // 0x0bbe
	13'h05e0: q3 = 16'h080b; // 0x0bc0
	13'h05e1: q3 = 16'h0c0d; // 0x0bc2
	13'h05e2: q3 = 16'h1010; // 0x0bc4
	13'h05e3: q3 = 16'h1010; // 0x0bc6
	13'h05e4: q3 = 16'h1010; // 0x0bc8
	13'h05e5: q3 = 16'h100d; // 0x0bca
	13'h05e6: q3 = 16'h0c0b; // 0x0bcc
	13'h05e7: q3 = 16'h0808; // 0x0bce
	13'h05e8: q3 = 16'h0001; // 0x0bd0
	13'h05e9: q3 = 16'h0000; // 0x0bd2
	13'h05ea: q3 = 16'h0000; // 0x0bd4
	13'h05eb: q3 = 16'h0007; // 0x0bd6
	13'h05ec: q3 = 16'h0608; // 0x0bd8
	13'h05ed: q3 = 16'h0706; // 0x0bda
	13'h05ee: q3 = 16'h0000; // 0x0bdc
	13'h05ef: q3 = 16'h0000; // 0x0bde
	13'h05f0: q3 = 16'h0000; // 0x0be0
	13'h05f1: q3 = 16'h0006; // 0x0be2
	13'h05f2: q3 = 16'h0708; // 0x0be4
	13'h05f3: q3 = 16'h0607; // 0x0be6
	13'h05f4: q3 = 16'h0000; // 0x0be8
	13'h05f5: q3 = 16'h0000; // 0x0bea
	13'h05f6: q3 = 16'h1313; // 0x0bec
	13'h05f7: q3 = 16'h1313; // 0x0bee
	13'h05f8: q3 = 16'h1313; // 0x0bf0
	13'h05f9: q3 = 16'h1313; // 0x0bf2
	13'h05fa: q3 = 16'h1211; // 0x0bf4
	13'h05fb: q3 = 16'h0f0d; // 0x0bf6
	13'h05fc: q3 = 16'h0b09; // 0x0bf8
	13'h05fd: q3 = 16'h0706; // 0x0bfa
	13'h05fe: q3 = 16'h0504; // 0x0bfc
	13'h05ff: q3 = 16'h0302; // 0x0bfe
	13'h0600: q3 = 16'h0100; // 0x0c00
	13'h0601: q3 = 16'h0000; // 0x0c02
	13'h0602: q3 = 16'h0102; // 0x0c04
	13'h0603: q3 = 16'h0304; // 0x0c06
	13'h0604: q3 = 16'h0506; // 0x0c08
	13'h0605: q3 = 16'h0708; // 0x0c0a
	13'h0606: q3 = 16'h0a0b; // 0x0c0c
	13'h0607: q3 = 16'h0b0b; // 0x0c0e
	13'h0608: q3 = 16'h0b0b; // 0x0c10
	13'h0609: q3 = 16'h0a08; // 0x0c12
	13'h060a: q3 = 16'h0706; // 0x0c14
	13'h060b: q3 = 16'h0504; // 0x0c16
	13'h060c: q3 = 16'h0302; // 0x0c18
	13'h060d: q3 = 16'h0100; // 0x0c1a
	13'h060e: q3 = 16'h0003; // 0x0c1c
	13'h060f: q3 = 16'h0004; // 0x0c1e
	13'h0610: q3 = 16'h0011; // 0x0c20
	13'h0611: q3 = 16'h0016; // 0x0c22
	13'h0612: q3 = 16'h0006; // 0x0c24
	13'h0613: q3 = 16'h0008; // 0x0c26
	13'h0614: q3 = 16'h000f; // 0x0c28
	13'h0615: q3 = 16'h0014; // 0x0c2a
	13'h0616: q3 = 16'h000d; // 0x0c2c
	13'h0617: q3 = 16'h000c; // 0x0c2e
	13'h0618: q3 = 16'h0506; // 0x0c30
	13'h0619: q3 = 16'h0707; // 0x0c32
	13'h061a: q3 = 16'h0708; // 0x0c34
	13'h061b: q3 = 16'h0808; // 0x0c36
	13'h061c: q3 = 16'h0707; // 0x0c38
	13'h061d: q3 = 16'h0606; // 0x0c3a
	13'h061e: q3 = 16'h0500; // 0x0c3c
	13'h061f: q3 = 16'h0303; // 0x0c3e
	13'h0620: q3 = 16'h0405; // 0x0c40
	13'h0621: q3 = 16'h0606; // 0x0c42
	13'h0622: q3 = 16'h0708; // 0x0c44
	13'h0623: q3 = 16'h0809; // 0x0c46
	13'h0624: q3 = 16'h090a; // 0x0c48
	13'h0625: q3 = 16'h0a00; // 0x0c4a
	13'h0626: q3 = 16'h0202; // 0x0c4c
	13'h0627: q3 = 16'h0102; // 0x0c4e
	13'h0628: q3 = 16'h0202; // 0x0c50
	13'h0629: q3 = 16'h0101; // 0x0c52
	13'h062a: q3 = 16'h0202; // 0x0c54
	13'h062b: q3 = 16'h0202; // 0x0c56
	13'h062c: q3 = 16'h0200; // 0x0c58
	13'h062d: q3 = 16'h0000; // 0x0c5a
	13'h062e: q3 = 16'h0001; // 0x0c5c
	13'h062f: q3 = 16'h0000; // 0x0c5e
	13'h0630: q3 = 16'h0000; // 0x0c60
	13'h0631: q3 = 16'h0000; // 0x0c62
	13'h0632: q3 = 16'h0000; // 0x0c64
	13'h0633: q3 = 16'h2020; // 0x0c66
	13'h0634: q3 = 16'h3000; // 0x0c68
	13'h0635: q3 = 16'h1416; // 0x0c6a
	13'h0636: q3 = 16'h1819; // 0x0c6c
	13'h0637: q3 = 16'h1a1a; // 0x0c6e
	13'h0638: q3 = 16'h1a1a; // 0x0c70
	13'h0639: q3 = 16'h1918; // 0x0c72
	13'h063a: q3 = 16'h1614; // 0x0c74
	13'h063b: q3 = 16'h110e; // 0x0c76
	13'h063c: q3 = 16'h0b09; // 0x0c78
	13'h063d: q3 = 16'h0706; // 0x0c7a
	13'h063e: q3 = 16'h0505; // 0x0c7c
	13'h063f: q3 = 16'h0505; // 0x0c7e
	13'h0640: q3 = 16'h0607; // 0x0c80
	13'h0641: q3 = 16'h090b; // 0x0c82
	13'h0642: q3 = 16'h0e11; // 0x0c84
	13'h0643: q3 = 16'h1c1b; // 0x0c86
	13'h0644: q3 = 16'h1a18; // 0x0c88
	13'h0645: q3 = 16'h1613; // 0x0c8a
	13'h0646: q3 = 16'h100d; // 0x0c8c
	13'h0647: q3 = 16'h0b09; // 0x0c8e
	13'h0648: q3 = 16'h0807; // 0x0c90
	13'h0649: q3 = 16'h0707; // 0x0c92
	13'h064a: q3 = 16'h0708; // 0x0c94
	13'h064b: q3 = 16'h090b; // 0x0c96
	13'h064c: q3 = 16'h0d10; // 0x0c98
	13'h064d: q3 = 16'h1316; // 0x0c9a
	13'h064e: q3 = 16'h181a; // 0x0c9c
	13'h064f: q3 = 16'h1b1c; // 0x0c9e
	13'h0650: q3 = 16'h1c1c; // 0x0ca0
	13'h0651: q3 = 16'h0000; // 0x0ca2
	13'h0652: q3 = 16'h0001; // 0x0ca4
	13'h0653: q3 = 16'h0000; // 0x0ca6
	13'h0654: q3 = 16'h0000; // 0x0ca8
	13'h0655: q3 = 16'h2000; // 0x0caa
	13'h0656: q3 = 16'h2000; // 0x0cac
	13'h0657: q3 = 16'h2100; // 0x0cae
	13'h0658: q3 = 16'h0909; // 0x0cb0
	13'h0659: q3 = 16'h0909; // 0x0cb2
	13'h065a: q3 = 16'h0909; // 0x0cb4
	13'h065b: q3 = 16'h0909; // 0x0cb6
	13'h065c: q3 = 16'h0909; // 0x0cb8
	13'h065d: q3 = 16'h0909; // 0x0cba
	13'h065e: q3 = 16'h0909; // 0x0cbc
	13'h065f: q3 = 16'h0909; // 0x0cbe
	13'h0660: q3 = 16'h0909; // 0x0cc0
	13'h0661: q3 = 16'h0909; // 0x0cc2
	13'h0662: q3 = 16'h0909; // 0x0cc4
	13'h0663: q3 = 16'h0909; // 0x0cc6
	13'h0664: q3 = 16'h0909; // 0x0cc8
	13'h0665: q3 = 16'h0909; // 0x0cca
	13'h0666: q3 = 16'h0909; // 0x0ccc
	13'h0667: q3 = 16'h0909; // 0x0cce
	13'h0668: q3 = 16'h0909; // 0x0cd0
	13'h0669: q3 = 16'h090b; // 0x0cd2
	13'h066a: q3 = 16'h2124; // 0x0cd4
	13'h066b: q3 = 16'h2424; // 0x0cd6
	13'h066c: q3 = 16'h2424; // 0x0cd8
	13'h066d: q3 = 16'h2424; // 0x0cda
	13'h066e: q3 = 16'h2424; // 0x0cdc
	13'h066f: q3 = 16'h2424; // 0x0cde
	13'h0670: q3 = 16'h2424; // 0x0ce0
	13'h0671: q3 = 16'h2424; // 0x0ce2
	13'h0672: q3 = 16'h2424; // 0x0ce4
	13'h0673: q3 = 16'h2424; // 0x0ce6
	13'h0674: q3 = 16'h2424; // 0x0ce8
	13'h0675: q3 = 16'h1715; // 0x0cea
	13'h0676: q3 = 16'h1515; // 0x0cec
	13'h0677: q3 = 16'h1515; // 0x0cee
	13'h0678: q3 = 16'h1516; // 0x0cf0
	13'h0679: q3 = 16'h181a; // 0x0cf2
	13'h067a: q3 = 16'h1a1b; // 0x0cf4
	13'h067b: q3 = 16'h1b1c; // 0x0cf6
	13'h067c: q3 = 16'h1d1e; // 0x0cf8
	13'h067d: q3 = 16'h1e1f; // 0x0cfa
	13'h067e: q3 = 16'h1f20; // 0x0cfc
	13'h067f: q3 = 16'h2122; // 0x0cfe
	13'h0680: q3 = 16'h2324; // 0x0d00
	13'h0681: q3 = 16'h2627; // 0x0d02
	13'h0682: q3 = 16'h2829; // 0x0d04
	13'h0683: q3 = 16'h2a2b; // 0x0d06
	13'h0684: q3 = 16'h2c2d; // 0x0d08
	13'h0685: q3 = 16'h2d2d; // 0x0d0a
	13'h0686: q3 = 16'h2e2e; // 0x0d0c
	13'h0687: q3 = 16'h2e30; // 0x0d0e
	13'h0688: q3 = 16'h3333; // 0x0d10
	13'h0689: q3 = 16'h3536; // 0x0d12
	13'h068a: q3 = 16'h3738; // 0x0d14
	13'h068b: q3 = 16'h393b; // 0x0d16
	13'h068c: q3 = 16'h3d3f; // 0x0d18
	13'h068d: q3 = 16'h3f3f; // 0x0d1a
	13'h068e: q3 = 16'h4041; // 0x0d1c
	13'h068f: q3 = 16'h4345; // 0x0d1e
	13'h0690: q3 = 16'h4600; // 0x0d20
	13'h0691: q3 = 16'h0001; // 0x0d22
	13'h0692: q3 = 16'h0203; // 0x0d24
	13'h0693: q3 = 16'h0303; // 0x0d26
	13'h0694: q3 = 16'h0303; // 0x0d28
	13'h0695: q3 = 16'h0303; // 0x0d2a
	13'h0696: q3 = 16'h0303; // 0x0d2c
	13'h0697: q3 = 16'h0303; // 0x0d2e
	13'h0698: q3 = 16'h0303; // 0x0d30
	13'h0699: q3 = 16'h0303; // 0x0d32
	13'h069a: q3 = 16'h0303; // 0x0d34
	13'h069b: q3 = 16'h0303; // 0x0d36
	13'h069c: q3 = 16'h0303; // 0x0d38
	13'h069d: q3 = 16'h0303; // 0x0d3a
	13'h069e: q3 = 16'h0303; // 0x0d3c
	13'h069f: q3 = 16'h0303; // 0x0d3e
	13'h06a0: q3 = 16'h0303; // 0x0d40
	13'h06a1: q3 = 16'h0303; // 0x0d42
	13'h06a2: q3 = 16'h0422; // 0x0d44
	13'h06a3: q3 = 16'h2525; // 0x0d46
	13'h06a4: q3 = 16'ha525; // 0x0d48
	13'h06a5: q3 = 16'h0504; // 0x0d4a
	13'h06a6: q3 = 16'h0404; // 0x0d4c
	13'h06a7: q3 = 16'h012e; // 0x0d4e
	13'h06a8: q3 = 16'haaaa; // 0x0d50
	13'h06a9: q3 = 16'h0000; // 0x0d52
	13'h06aa: q3 = 16'h0000; // 0x0d54
	13'h06ab: q3 = 16'h26a7; // 0x0d56
	13'h06ac: q3 = 16'h2728; // 0x0d58
	13'h06ad: q3 = 16'h0000; // 0x0d5a
	13'h06ae: q3 = 16'h2524; // 0x0d5c
	13'h06af: q3 = 16'h2324; // 0x0d5e
	13'h06b0: q3 = 16'h2424; // 0x0d60
	13'h06b1: q3 = 16'h24a4; // 0x0d62
	13'h06b2: q3 = 16'ha426; // 0x0d64
	13'h06b3: q3 = 16'h393e; // 0x0d66
	13'h06b4: q3 = 16'h3e3e; // 0x0d68
	13'h06b5: q3 = 16'h3e3e; // 0x0d6a
	13'h06b6: q3 = 16'h3e3c; // 0x0d6c
	13'h06b7: q3 = 16'h3b3a; // 0x0d6e
	13'h06b8: q3 = 16'h3a3a; // 0x0d70
	13'h06b9: q3 = 16'h3a3a; // 0x0d72
	13'h06ba: q3 = 16'h3a3a; // 0x0d74
	13'h06bb: q3 = 16'h3a3a; // 0x0d76
	13'h06bc: q3 = 16'h3b3a; // 0x0d78
	13'h06bd: q3 = 16'h3a3a; // 0x0d7a
	13'h06be: q3 = 16'h3939; // 0x0d7c
	13'h06bf: q3 = 16'h3939; // 0x0d7e
	13'h06c0: q3 = 16'h3635; // 0x0d80
	13'h06c1: q3 = 16'h32ae; // 0x0d82
	13'h06c2: q3 = 16'habaa; // 0x0d84
	13'h06c3: q3 = 16'ha8a7; // 0x0d86
	13'h06c4: q3 = 16'ha4a1; // 0x0d88
	13'h06c5: q3 = 16'ha09d; // 0x0d8a
	13'h06c6: q3 = 16'h9c9b; // 0x0d8c
	13'h06c7: q3 = 16'h9999; // 0x0d8e
	13'h06c8: q3 = 16'h9795; // 0x0d90
	13'h06c9: q3 = 16'h9292; // 0x0d92
	13'h06ca: q3 = 16'h9292; // 0x0d94
	13'h06cb: q3 = 16'h9599; // 0x0d96
	13'h06cc: q3 = 16'h9da2; // 0x0d98
	13'h06cd: q3 = 16'ha5a9; // 0x0d9a
	13'h06ce: q3 = 16'habac; // 0x0d9c
	13'h06cf: q3 = 16'haba4; // 0x0d9e
	13'h06d0: q3 = 16'h9c9a; // 0x0da0
	13'h06d1: q3 = 16'h1a1c; // 0x0da2
	13'h06d2: q3 = 16'h1f20; // 0x0da4
	13'h06d3: q3 = 16'h2020; // 0x0da6
	13'h06d4: q3 = 16'h2020; // 0x0da8
	13'h06d5: q3 = 16'h2020; // 0x0daa
	13'h06d6: q3 = 16'h2020; // 0x0dac
	13'h06d7: q3 = 16'h2020; // 0x0dae
	13'h06d8: q3 = 16'h2020; // 0x0db0
	13'h06d9: q3 = 16'h2021; // 0x0db2
	13'h06da: q3 = 16'h2121; // 0x0db4
	13'h06db: q3 = 16'h2121; // 0x0db6
	13'h06dc: q3 = 16'h2121; // 0x0db8
	13'h06dd: q3 = 16'h2121; // 0x0dba
	13'h06de: q3 = 16'h2121; // 0x0dbc
	13'h06df: q3 = 16'h2121; // 0x0dbe
	13'h06e0: q3 = 16'h2121; // 0x0dc0
	13'h06e1: q3 = 16'h2121; // 0x0dc2
	13'h06e2: q3 = 16'h2121; // 0x0dc4
	13'h06e3: q3 = 16'h2121; // 0x0dc6
	13'h06e4: q3 = 16'h0b03; // 0x0dc8
	13'h06e5: q3 = 16'h0404; // 0x0dca
	13'h06e6: q3 = 16'h0403; // 0x0dcc
	13'h06e7: q3 = 16'h0304; // 0x0dce
	13'h06e8: q3 = 16'h0403; // 0x0dd0
	13'h06e9: q3 = 16'h0303; // 0x0dd2
	13'h06ea: q3 = 16'h0304; // 0x0dd4
	13'h06eb: q3 = 16'h0507; // 0x0dd6
	13'h06ec: q3 = 16'h0707; // 0x0dd8
	13'h06ed: q3 = 16'h0808; // 0x0dda
	13'h06ee: q3 = 16'h0809; // 0x0ddc
	13'h06ef: q3 = 16'h0909; // 0x0dde
	13'h06f0: q3 = 16'h090a; // 0x0de0
	13'h06f1: q3 = 16'h0c0d; // 0x0de2
	13'h06f2: q3 = 16'h0d0d; // 0x0de4
	13'h06f3: q3 = 16'h0e10; // 0x0de6
	13'h06f4: q3 = 16'h1316; // 0x0de8
	13'h06f5: q3 = 16'h191b; // 0x0dea
	13'h06f6: q3 = 16'h1b1b; // 0x0dec
	13'h06f7: q3 = 16'h1b1b; // 0x0dee
	13'h06f8: q3 = 16'h1b1b; // 0x0df0
	13'h06f9: q3 = 16'h1b1b; // 0x0df2
	13'h06fa: q3 = 16'h1b1b; // 0x0df4
	13'h06fb: q3 = 16'h1b1d; // 0x0df6
	13'h06fc: q3 = 16'h1d1f; // 0x0df8
	13'h06fd: q3 = 16'h2124; // 0x0dfa
	13'h06fe: q3 = 16'h2627; // 0x0dfc
	13'h06ff: q3 = 16'h292b; // 0x0dfe
	13'h0700: q3 = 16'h2c2c; // 0x0e00
	13'h0701: q3 = 16'h2c2c; // 0x0e02
	13'h0702: q3 = 16'h2c2c; // 0x0e04
	13'h0703: q3 = 16'h2c2c; // 0x0e06
	13'h0704: q3 = 16'h2c2c; // 0x0e08
	13'h0705: q3 = 16'h2d2d; // 0x0e0a
	13'h0706: q3 = 16'h2e30; // 0x0e0c
	13'h0707: q3 = 16'h3233; // 0x0e0e
	13'h0708: q3 = 16'h3333; // 0x0e10
	13'h0709: q3 = 16'h3333; // 0x0e12
	13'h070a: q3 = 16'h3333; // 0x0e14
	13'h070b: q3 = 16'h3333; // 0x0e16
	13'h070c: q3 = 16'h3333; // 0x0e18
	13'h070d: q3 = 16'h3333; // 0x0e1a
	13'h070e: q3 = 16'h3333; // 0x0e1c
	13'h070f: q3 = 16'h3230; // 0x0e1e
	13'h0710: q3 = 16'h302e; // 0x0e20
	13'h0711: q3 = 16'h2d2d; // 0x0e22
	13'h0712: q3 = 16'h2d2c; // 0x0e24
	13'h0713: q3 = 16'h2a27; // 0x0e26
	13'h0714: q3 = 16'h2421; // 0x0e28
	13'h0715: q3 = 16'h9a19; // 0x0e2a
	13'h0716: q3 = 16'h1919; // 0x0e2c
	13'h0717: q3 = 16'h1919; // 0x0e2e
	13'h0718: q3 = 16'h1919; // 0x0e30
	13'h0719: q3 = 16'h1919; // 0x0e32
	13'h071a: q3 = 16'h1919; // 0x0e34
	13'h071b: q3 = 16'h1919; // 0x0e36
	13'h071c: q3 = 16'h1900; // 0x0e38
	13'h071d: q3 = 16'hffff; // 0x0e3a
	13'h071e: q3 = 16'hffff; // 0x0e3c
	13'h071f: q3 = 16'hffff; // 0x0e3e
	13'h0720: q3 = 16'hffff; // 0x0e40
	13'h0721: q3 = 16'hffff; // 0x0e42
	13'h0722: q3 = 16'hffff; // 0x0e44
	13'h0723: q3 = 16'hffff; // 0x0e46
	13'h0724: q3 = 16'hffff; // 0x0e48
	13'h0725: q3 = 16'hffff; // 0x0e4a
	13'h0726: q3 = 16'hfcb7; // 0x0e4c
	13'h0727: q3 = 16'hfd1e; // 0x0e4e
	13'h0728: q3 = 16'hf9ff; // 0x0e50
	13'h0729: q3 = 16'hffff; // 0x0e52
	13'h072a: q3 = 16'h3000; // 0x0e54
	13'h072b: q3 = 16'h0000; // 0x0e56
	13'h072c: q3 = 16'h0fff; // 0x0e58
	13'h072d: q3 = 16'hffff; // 0x0e5a
	13'h072e: q3 = 16'h7ffe; // 0x0e5c
	13'h072f: q3 = 16'hffff; // 0x0e5e
	13'h0730: q3 = 16'hffff; // 0x0e60
	13'h0731: q3 = 16'hffff; // 0x0e62
	13'h0732: q3 = 16'hffff; // 0x0e64
	13'h0733: q3 = 16'hffff; // 0x0e66
	13'h0734: q3 = 16'hffff; // 0x0e68
	13'h0735: q3 = 16'hffff; // 0x0e6a
	13'h0736: q3 = 16'h0000; // 0x0e6c
	13'h0737: q3 = 16'h0078; // 0x0e6e
	13'h0738: q3 = 16'h0000; // 0x0e70
	13'h0739: q3 = 16'h0000; // 0x0e72
	13'h073a: q3 = 16'h0000; // 0x0e74
	13'h073b: q3 = 16'h6dc6; // 0x0e76
	13'h073c: q3 = 16'h0000; // 0x0e78
	13'h073d: q3 = 16'h6de8; // 0x0e7a
	13'h073e: q3 = 16'h0000; // 0x0e7c
	13'h073f: q3 = 16'h6e08; // 0x0e7e
	13'h0740: q3 = 16'h0000; // 0x0e80
	13'h0741: q3 = 16'h6e28; // 0x0e82
	13'h0742: q3 = 16'h4f53; // 0x0e84
	13'h0743: q3 = 16'h4341; // 0x0e86
	13'h0744: q3 = 16'h5200; // 0x0e88
	13'h0745: q3 = 16'h414e; // 0x0e8a
	13'h0746: q3 = 16'h4745; // 0x0e8c
	13'h0747: q3 = 16'h4c4f; // 0x0e8e
	13'h0748: q3 = 16'h004a; // 0x0e90
	13'h0749: q3 = 16'h4143; // 0x0e92
	13'h074a: q3 = 16'h5155; // 0x0e94
	13'h074b: q3 = 16'h4553; // 0x0e96
	13'h074c: q3 = 16'h005a; // 0x0e98
	13'h074d: q3 = 16'h4f52; // 0x0e9a
	13'h074e: q3 = 16'h4241; // 0x0e9c
	13'h074f: q3 = 16'h0020; // 0x0e9e
	13'h0750: q3 = 16'h2020; // 0x0ea0
	13'h0751: q3 = 16'h2043; // 0x0ea2
	13'h0752: q3 = 16'h4841; // 0x0ea4
	13'h0753: q3 = 16'h524c; // 0x0ea6
	13'h0754: q3 = 16'h4559; // 0x0ea8
	13'h0755: q3 = 16'h2043; // 0x0eaa
	13'h0756: q3 = 16'h4855; // 0x0eac
	13'h0757: q3 = 16'h434b; // 0x0eae
	13'h0758: q3 = 16'h2020; // 0x0eb0
	13'h0759: q3 = 16'h0050; // 0x0eb2
	13'h075a: q3 = 16'h4f55; // 0x0eb4
	13'h075b: q3 = 16'h5200; // 0x0eb6
	13'h075c: q3 = 16'h0095; // 0x0eb8
	13'h075d: q3 = 16'h8000; // 0x0eba
	13'h075e: q3 = 16'h0094; // 0x0ebc
	13'h075f: q3 = 16'h8000; // 0x0ebe
	13'h0760: q3 = 16'h00a8; // 0x0ec0
	13'h0761: q3 = 16'h0000; // 0x0ec2
	13'h0762: q3 = 16'h0094; // 0x0ec4
	13'h0763: q3 = 16'h0000; // 0x0ec6
	13'h0764: q3 = 16'h0094; // 0x0ec8
	13'h0765: q3 = 16'h4000; // 0x0eca
	13'h0766: q3 = 16'h0094; // 0x0ecc
	13'h0767: q3 = 16'h4004; // 0x0ece
	13'h0768: q3 = 16'h0094; // 0x0ed0
	13'h0769: q3 = 16'h4002; // 0x0ed2
	13'h076a: q3 = 16'h0094; // 0x0ed4
	13'h076b: q3 = 16'h4006; // 0x0ed6
	13'h076c: q3 = 16'h0094; // 0x0ed8
	13'h076d: q3 = 16'hc000; // 0x0eda
	13'h076e: q3 = 16'h000f; // 0x0edc
	13'h076f: q3 = 16'h0200; // 0x0ede
	13'h0770: q3 = 16'h003a; // 0x0ee0
	13'h0771: q3 = 16'haaaa; // 0x0ee2
	13'h0772: q3 = 16'h030f; // 0x0ee4
	13'h0773: q3 = 16'h0000; // 0x0ee6
	13'h0774: q3 = 16'hf332; // 0x0ee8
	13'h0775: q3 = 16'h0000; // 0x0eea
	13'h0776: q3 = 16'hc314; // 0x0eec
	13'h0777: q3 = 16'h0000; // 0x0eee
	13'h0778: q3 = 16'hc338; // 0x0ef0
	13'h0779: q3 = 16'h0000; // 0x0ef2
	13'h077a: q3 = 16'hc338; // 0x0ef4
	13'h077b: q3 = 16'h050f; // 0x0ef6
	13'h077c: q3 = 16'h0000; // 0x0ef8
	13'h077d: q3 = 16'hf34a; // 0x0efa
	13'h077e: q3 = 16'h0000; // 0x0efc
	13'h077f: q3 = 16'hc320; // 0x0efe
	13'h0780: q3 = 16'h0000; // 0x0f00
	13'h0781: q3 = 16'hc350; // 0x0f02
	13'h0782: q3 = 16'h0000; // 0x0f04
	13'h0783: q3 = 16'hc350; // 0x0f06
	13'h0784: q3 = 16'h0d00; // 0x0f08
	13'h0785: q3 = 16'h0000; // 0x0f0a
	13'h0786: q3 = 16'hd4b0; // 0x0f0c
	13'h0787: q3 = 16'h080f; // 0x0f0e
	13'h0788: q3 = 16'h0100; // 0x0f10
	13'h0789: q3 = 16'h0005; // 0x0f12
	13'h078a: q3 = 16'h0d01; // 0x0f14
	13'h078b: q3 = 16'h0000; // 0x0f16
	13'h078c: q3 = 16'hd0e8; // 0x0f18
	13'h078d: q3 = 16'h0002; // 0x0f1a
	13'h078e: q3 = 16'h0d01; // 0x0f1c
	13'h078f: q3 = 16'h0000; // 0x0f1e
	13'h0790: q3 = 16'hd1da; // 0x0f20
	13'h0791: q3 = 16'h0d01; // 0x0f22
	13'h0792: q3 = 16'h0000; // 0x0f24
	13'h0793: q3 = 16'hd76a; // 0x0f26
	13'h0794: q3 = 16'h0d00; // 0x0f28
	13'h0795: q3 = 16'h0000; // 0x0f2a
	13'h0796: q3 = 16'hd1da; // 0x0f2c
	13'h0797: q3 = 16'h0d00; // 0x0f2e
	13'h0798: q3 = 16'h0000; // 0x0f30
	13'h0799: q3 = 16'hd874; // 0x0f32
	13'h079a: q3 = 16'h0008; // 0x0f34
	13'h079b: q3 = 16'h0d00; // 0x0f36
	13'h079c: q3 = 16'h0000; // 0x0f38
	13'h079d: q3 = 16'hd4b0; // 0x0f3a
	13'h079e: q3 = 16'h080f; // 0x0f3c
	13'h079f: q3 = 16'h0100; // 0x0f3e
	13'h07a0: q3 = 16'h0005; // 0x0f40
	13'h07a1: q3 = 16'h0d01; // 0x0f42
	13'h07a2: q3 = 16'h0000; // 0x0f44
	13'h07a3: q3 = 16'hd0e8; // 0x0f46
	13'h07a4: q3 = 16'h0002; // 0x0f48
	13'h07a5: q3 = 16'h0d01; // 0x0f4a
	13'h07a6: q3 = 16'h0000; // 0x0f4c
	13'h07a7: q3 = 16'hd1da; // 0x0f4e
	13'h07a8: q3 = 16'h0d01; // 0x0f50
	13'h07a9: q3 = 16'h0000; // 0x0f52
	13'h07aa: q3 = 16'hd76a; // 0x0f54
	13'h07ab: q3 = 16'h0008; // 0x0f56
	13'h07ac: q3 = 16'h0d00; // 0x0f58
	13'h07ad: q3 = 16'h0000; // 0x0f5a
	13'h07ae: q3 = 16'hd64a; // 0x0f5c
	13'h07af: q3 = 16'h0d00; // 0x0f5e
	13'h07b0: q3 = 16'h0000; // 0x0f60
	13'h07b1: q3 = 16'hd2dc; // 0x0f62
	13'h07b2: q3 = 16'h0d00; // 0x0f64
	13'h07b3: q3 = 16'h0000; // 0x0f66
	13'h07b4: q3 = 16'hd58c; // 0x0f68
	13'h07b5: q3 = 16'h0d00; // 0x0f6a
	13'h07b6: q3 = 16'h0000; // 0x0f6c
	13'h07b7: q3 = 16'hd4b0; // 0x0f6e
	13'h07b8: q3 = 16'h080f; // 0x0f70
	13'h07b9: q3 = 16'h0100; // 0x0f72
	13'h07ba: q3 = 16'h0005; // 0x0f74
	13'h07bb: q3 = 16'h0d01; // 0x0f76
	13'h07bc: q3 = 16'h0000; // 0x0f78
	13'h07bd: q3 = 16'hd0e8; // 0x0f7a
	13'h07be: q3 = 16'h0002; // 0x0f7c
	13'h07bf: q3 = 16'h0d01; // 0x0f7e
	13'h07c0: q3 = 16'h0000; // 0x0f80
	13'h07c1: q3 = 16'hd1da; // 0x0f82
	13'h07c2: q3 = 16'h0d00; // 0x0f84
	13'h07c3: q3 = 16'h0000; // 0x0f86
	13'h07c4: q3 = 16'hd874; // 0x0f88
	13'h07c5: q3 = 16'h0d00; // 0x0f8a
	13'h07c6: q3 = 16'h0000; // 0x0f8c
	13'h07c7: q3 = 16'hd904; // 0x0f8e
	13'h07c8: q3 = 16'h0008; // 0x0f90
	13'h07c9: q3 = 16'h0d00; // 0x0f92
	13'h07ca: q3 = 16'h0000; // 0x0f94
	13'h07cb: q3 = 16'hd96e; // 0x0f96
	13'h07cc: q3 = 16'h0d00; // 0x0f98
	13'h07cd: q3 = 16'h0000; // 0x0f9a
	13'h07ce: q3 = 16'hd4b0; // 0x0f9c
	13'h07cf: q3 = 16'h080f; // 0x0f9e
	13'h07d0: q3 = 16'h0100; // 0x0fa0
	13'h07d1: q3 = 16'h0005; // 0x0fa2
	13'h07d2: q3 = 16'h0d01; // 0x0fa4
	13'h07d3: q3 = 16'h0000; // 0x0fa6
	13'h07d4: q3 = 16'hd0e8; // 0x0fa8
	13'h07d5: q3 = 16'h0002; // 0x0faa
	13'h07d6: q3 = 16'h0d01; // 0x0fac
	13'h07d7: q3 = 16'h0000; // 0x0fae
	13'h07d8: q3 = 16'hd1da; // 0x0fb0
	13'h07d9: q3 = 16'h0d01; // 0x0fb2
	13'h07da: q3 = 16'h0000; // 0x0fb4
	13'h07db: q3 = 16'hd76a; // 0x0fb6
	13'h07dc: q3 = 16'h0d00; // 0x0fb8
	13'h07dd: q3 = 16'h0000; // 0x0fba
	13'h07de: q3 = 16'hd1da; // 0x0fbc
	13'h07df: q3 = 16'h0d00; // 0x0fbe
	13'h07e0: q3 = 16'h0000; // 0x0fc0
	13'h07e1: q3 = 16'hd874; // 0x0fc2
	13'h07e2: q3 = 16'h0d00; // 0x0fc4
	13'h07e3: q3 = 16'h0000; // 0x0fc6
	13'h07e4: q3 = 16'hd904; // 0x0fc8
	13'h07e5: q3 = 16'h0008; // 0x0fca
	13'h07e6: q3 = 16'h0d00; // 0x0fcc
	13'h07e7: q3 = 16'h0000; // 0x0fce
	13'h07e8: q3 = 16'hd64a; // 0x0fd0
	13'h07e9: q3 = 16'h0d00; // 0x0fd2
	13'h07ea: q3 = 16'h0000; // 0x0fd4
	13'h07eb: q3 = 16'hd2dc; // 0x0fd6
	13'h07ec: q3 = 16'h0d00; // 0x0fd8
	13'h07ed: q3 = 16'h0000; // 0x0fda
	13'h07ee: q3 = 16'hd64a; // 0x0fdc
	13'h07ef: q3 = 16'h0d00; // 0x0fde
	13'h07f0: q3 = 16'h0000; // 0x0fe0
	13'h07f1: q3 = 16'hd410; // 0x0fe2
	13'h07f2: q3 = 16'h0d00; // 0x0fe4
	13'h07f3: q3 = 16'h0000; // 0x0fe6
	13'h07f4: q3 = 16'hd4b0; // 0x0fe8
	13'h07f5: q3 = 16'h080f; // 0x0fea
	13'h07f6: q3 = 16'h0100; // 0x0fec
	13'h07f7: q3 = 16'h0005; // 0x0fee
	13'h07f8: q3 = 16'h0d01; // 0x0ff0
	13'h07f9: q3 = 16'h0000; // 0x0ff2
	13'h07fa: q3 = 16'hd0e8; // 0x0ff4
	13'h07fb: q3 = 16'h0002; // 0x0ff6
	13'h07fc: q3 = 16'h0d01; // 0x0ff8
	13'h07fd: q3 = 16'h0000; // 0x0ffa
	13'h07fe: q3 = 16'hd1da; // 0x0ffc
	13'h07ff: q3 = 16'h0d01; // 0x0ffe
	13'h0800: q3 = 16'h0000; // 0x1000
	13'h0801: q3 = 16'hd76a; // 0x1002
	13'h0802: q3 = 16'h0d00; // 0x1004
	13'h0803: q3 = 16'h0000; // 0x1006
	13'h0804: q3 = 16'hd1da; // 0x1008
	13'h0805: q3 = 16'h0d00; // 0x100a
	13'h0806: q3 = 16'h0000; // 0x100c
	13'h0807: q3 = 16'hd874; // 0x100e
	13'h0808: q3 = 16'h0d00; // 0x1010
	13'h0809: q3 = 16'h0000; // 0x1012
	13'h080a: q3 = 16'hd904; // 0x1014
	13'h080b: q3 = 16'h0008; // 0x1016
	13'h080c: q3 = 16'h0d00; // 0x1018
	13'h080d: q3 = 16'h0000; // 0x101a
	13'h080e: q3 = 16'hd96e; // 0x101c
	13'h080f: q3 = 16'h0d00; // 0x101e
	13'h0810: q3 = 16'h0000; // 0x1020
	13'h0811: q3 = 16'hd61e; // 0x1022
	13'h0812: q3 = 16'h0d00; // 0x1024
	13'h0813: q3 = 16'h0000; // 0x1026
	13'h0814: q3 = 16'hd4b0; // 0x1028
	13'h0815: q3 = 16'h080f; // 0x102a
	13'h0816: q3 = 16'h0100; // 0x102c
	13'h0817: q3 = 16'h0005; // 0x102e
	13'h0818: q3 = 16'h0d01; // 0x1030
	13'h0819: q3 = 16'h0000; // 0x1032
	13'h081a: q3 = 16'hd0e8; // 0x1034
	13'h081b: q3 = 16'h0002; // 0x1036
	13'h081c: q3 = 16'h0d01; // 0x1038
	13'h081d: q3 = 16'h0000; // 0x103a
	13'h081e: q3 = 16'hd1da; // 0x103c
	13'h081f: q3 = 16'h0d00; // 0x103e
	13'h0820: q3 = 16'h0000; // 0x1040
	13'h0821: q3 = 16'hd874; // 0x1042
	13'h0822: q3 = 16'h0d00; // 0x1044
	13'h0823: q3 = 16'h0000; // 0x1046
	13'h0824: q3 = 16'hd904; // 0x1048
	13'h0825: q3 = 16'h0008; // 0x104a
	13'h0826: q3 = 16'h0d00; // 0x104c
	13'h0827: q3 = 16'h0000; // 0x104e
	13'h0828: q3 = 16'hd96e; // 0x1050
	13'h0829: q3 = 16'h0d00; // 0x1052
	13'h082a: q3 = 16'h0000; // 0x1054
	13'h082b: q3 = 16'hd64a; // 0x1056
	13'h082c: q3 = 16'h0d00; // 0x1058
	13'h082d: q3 = 16'h0000; // 0x105a
	13'h082e: q3 = 16'hd2dc; // 0x105c
	13'h082f: q3 = 16'h0d00; // 0x105e
	13'h0830: q3 = 16'h0000; // 0x1060
	13'h0831: q3 = 16'hd64a; // 0x1062
	13'h0832: q3 = 16'h0d00; // 0x1064
	13'h0833: q3 = 16'h0000; // 0x1066
	13'h0834: q3 = 16'hd410; // 0x1068
	13'h0835: q3 = 16'h0d00; // 0x106a
	13'h0836: q3 = 16'h0000; // 0x106c
	13'h0837: q3 = 16'hd4b0; // 0x106e
	13'h0838: q3 = 16'h080f; // 0x1070
	13'h0839: q3 = 16'h0100; // 0x1072
	13'h083a: q3 = 16'h0005; // 0x1074
	13'h083b: q3 = 16'h0d01; // 0x1076
	13'h083c: q3 = 16'h0000; // 0x1078
	13'h083d: q3 = 16'hd0e8; // 0x107a
	13'h083e: q3 = 16'h0002; // 0x107c
	13'h083f: q3 = 16'h0d01; // 0x107e
	13'h0840: q3 = 16'h0000; // 0x1080
	13'h0841: q3 = 16'hd1da; // 0x1082
	13'h0842: q3 = 16'h0d00; // 0x1084
	13'h0843: q3 = 16'h0000; // 0x1086
	13'h0844: q3 = 16'hd76a; // 0x1088
	13'h0845: q3 = 16'h0d00; // 0x108a
	13'h0846: q3 = 16'h0000; // 0x108c
	13'h0847: q3 = 16'hd58c; // 0x108e
	13'h0848: q3 = 16'h0d00; // 0x1090
	13'h0849: q3 = 16'h0000; // 0x1092
	13'h084a: q3 = 16'hd904; // 0x1094
	13'h084b: q3 = 16'h0008; // 0x1096
	13'h084c: q3 = 16'h0d00; // 0x1098
	13'h084d: q3 = 16'h0000; // 0x109a
	13'h084e: q3 = 16'hd96e; // 0x109c
	13'h084f: q3 = 16'h0d00; // 0x109e
	13'h0850: q3 = 16'h0000; // 0x10a0
	13'h0851: q3 = 16'hd64a; // 0x10a2
	13'h0852: q3 = 16'h0d00; // 0x10a4
	13'h0853: q3 = 16'h0000; // 0x10a6
	13'h0854: q3 = 16'hd2dc; // 0x10a8
	13'h0855: q3 = 16'h0d00; // 0x10aa
	13'h0856: q3 = 16'h0000; // 0x10ac
	13'h0857: q3 = 16'hd64a; // 0x10ae
	13'h0858: q3 = 16'h0d00; // 0x10b0
	13'h0859: q3 = 16'h0000; // 0x10b2
	13'h085a: q3 = 16'hd410; // 0x10b4
	13'h085b: q3 = 16'h0d00; // 0x10b6
	13'h085c: q3 = 16'h0000; // 0x10b8
	13'h085d: q3 = 16'hd4b0; // 0x10ba
	13'h085e: q3 = 16'h080f; // 0x10bc
	13'h085f: q3 = 16'h0100; // 0x10be
	13'h0860: q3 = 16'h0005; // 0x10c0
	13'h0861: q3 = 16'h0d01; // 0x10c2
	13'h0862: q3 = 16'h0000; // 0x10c4
	13'h0863: q3 = 16'hd0e8; // 0x10c6
	13'h0864: q3 = 16'h0002; // 0x10c8
	13'h0865: q3 = 16'h0d01; // 0x10ca
	13'h0866: q3 = 16'h0000; // 0x10cc
	13'h0867: q3 = 16'hd1da; // 0x10ce
	13'h0868: q3 = 16'h0d01; // 0x10d0
	13'h0869: q3 = 16'h0000; // 0x10d2
	13'h086a: q3 = 16'hd76a; // 0x10d4
	13'h086b: q3 = 16'h0d00; // 0x10d6
	13'h086c: q3 = 16'h0000; // 0x10d8
	13'h086d: q3 = 16'hd58c; // 0x10da
	13'h086e: q3 = 16'h0008; // 0x10dc
	13'h086f: q3 = 16'h0d00; // 0x10de
	13'h0870: q3 = 16'h0000; // 0x10e0
	13'h0871: q3 = 16'hd4b0; // 0x10e2
	13'h0872: q3 = 16'h080f; // 0x10e4
	13'h0873: q3 = 16'h0100; // 0x10e6
	13'h0874: q3 = 16'h030f; // 0x10e8
	13'h0875: q3 = 16'h0000; // 0x10ea
	13'h0876: q3 = 16'hf332; // 0x10ec
	13'h0877: q3 = 16'h0000; // 0x10ee
	13'h0878: q3 = 16'hc314; // 0x10f0
	13'h0879: q3 = 16'h0000; // 0x10f2
	13'h087a: q3 = 16'hc338; // 0x10f4
	13'h087b: q3 = 16'h0000; // 0x10f6
	13'h087c: q3 = 16'hc338; // 0x10f8
	13'h087d: q3 = 16'h050f; // 0x10fa
	13'h087e: q3 = 16'h0000; // 0x10fc
	13'h087f: q3 = 16'hf34a; // 0x10fe
	13'h0880: q3 = 16'h0000; // 0x1100
	13'h0881: q3 = 16'hc320; // 0x1102
	13'h0882: q3 = 16'h0000; // 0x1104
	13'h0883: q3 = 16'hc350; // 0x1106
	13'h0884: q3 = 16'h0000; // 0x1108
	13'h0885: q3 = 16'hc350; // 0x110a
	13'h0886: q3 = 16'h8705; // 0x110c
	13'h0887: q3 = 16'h0199; // 0x110e
	13'h0888: q3 = 16'h0333; // 0x1110
	13'h0889: q3 = 16'h0400; // 0x1112
	13'h088a: q3 = 16'h8b01; // 0x1114
	13'h088b: q3 = 16'h01b1; // 0x1116
	13'h088c: q3 = 16'h0400; // 0x1118
	13'h088d: q3 = 16'h8701; // 0x111a
	13'h088e: q3 = 16'h0199; // 0x111c
	13'h088f: q3 = 16'h0400; // 0x111e
	13'h0890: q3 = 16'h8701; // 0x1120
	13'h0891: q3 = 16'h0145; // 0x1122
	13'h0892: q3 = 16'h0400; // 0x1124
	13'h0893: q3 = 16'h8705; // 0x1126
	13'h0894: q3 = 16'h0222; // 0x1128
	13'h0895: q3 = 16'h0445; // 0x112a
	13'h0896: q3 = 16'h0400; // 0x112c
	13'h0897: q3 = 16'h8b01; // 0x112e
	13'h0898: q3 = 16'h0243; // 0x1130
	13'h0899: q3 = 16'h0400; // 0x1132
	13'h089a: q3 = 16'h8701; // 0x1134
	13'h089b: q3 = 16'h0222; // 0x1136
	13'h089c: q3 = 16'h0400; // 0x1138
	13'h089d: q3 = 16'h8701; // 0x113a
	13'h089e: q3 = 16'h0199; // 0x113c
	13'h089f: q3 = 16'h0400; // 0x113e
	13'h08a0: q3 = 16'h8705; // 0x1140
	13'h08a1: q3 = 16'h028a; // 0x1142
	13'h08a2: q3 = 16'h0514; // 0x1144
	13'h08a3: q3 = 16'h0400; // 0x1146
	13'h08a4: q3 = 16'h8b01; // 0x1148
	13'h08a5: q3 = 16'h02b0; // 0x114a
	13'h08a6: q3 = 16'h0400; // 0x114c
	13'h08a7: q3 = 16'h8701; // 0x114e
	13'h08a8: q3 = 16'h028a; // 0x1150
	13'h08a9: q3 = 16'h0400; // 0x1152
	13'h08aa: q3 = 16'h8701; // 0x1154
	13'h08ab: q3 = 16'h0222; // 0x1156
	13'h08ac: q3 = 16'h0400; // 0x1158
	13'h08ad: q3 = 16'h8705; // 0x115a
	13'h08ae: q3 = 16'h0333; // 0x115c
	13'h08af: q3 = 16'h0666; // 0x115e
	13'h08b0: q3 = 16'h0400; // 0x1160
	13'h08b1: q3 = 16'h8b01; // 0x1162
	13'h08b2: q3 = 16'h0363; // 0x1164
	13'h08b3: q3 = 16'h0400; // 0x1166
	13'h08b4: q3 = 16'h8701; // 0x1168
	13'h08b5: q3 = 16'h0333; // 0x116a
	13'h08b6: q3 = 16'h0400; // 0x116c
	13'h08b7: q3 = 16'h8701; // 0x116e
	13'h08b8: q3 = 16'h028a; // 0x1170
	13'h08b9: q3 = 16'h0400; // 0x1172
	13'h08ba: q3 = 16'h8705; // 0x1174
	13'h08bb: q3 = 16'h0445; // 0x1176
	13'h08bc: q3 = 16'h088b; // 0x1178
	13'h08bd: q3 = 16'h0900; // 0x117a
	13'h08be: q3 = 16'h8a05; // 0x117c
	13'h08bf: q3 = 16'h0300; // 0x117e
	13'h08c0: q3 = 16'h8705; // 0x1180
	13'h08c1: q3 = 16'h0408; // 0x1182
	13'h08c2: q3 = 16'h0810; // 0x1184
	13'h08c3: q3 = 16'h0300; // 0x1186
	13'h08c4: q3 = 16'h8a05; // 0x1188
	13'h08c5: q3 = 16'h0100; // 0x118a
	13'h08c6: q3 = 16'h8705; // 0x118c
	13'h08c7: q3 = 16'h03ce; // 0x118e
	13'h08c8: q3 = 16'h079c; // 0x1190
	13'h08c9: q3 = 16'h0400; // 0x1192
	13'h08ca: q3 = 16'h8a05; // 0x1194
	13'h08cb: q3 = 16'h0400; // 0x1196
	13'h08cc: q3 = 16'h8705; // 0x1198
	13'h08cd: q3 = 16'h0397; // 0x119a
	13'h08ce: q3 = 16'h072f; // 0x119c
	13'h08cf: q3 = 16'h0400; // 0x119e
	13'h08d0: q3 = 16'h8a05; // 0x11a0
	13'h08d1: q3 = 16'h0400; // 0x11a2
	13'h08d2: q3 = 16'h8705; // 0x11a4
	13'h08d3: q3 = 16'h0363; // 0x11a6
	13'h08d4: q3 = 16'h06c7; // 0x11a8
	13'h08d5: q3 = 16'h0800; // 0x11aa
	13'h08d6: q3 = 16'h8a04; // 0x11ac
	13'h08d7: q3 = 16'h0400; // 0x11ae
	13'h08d8: q3 = 16'h0601; // 0x11b0
	13'h08d9: q3 = 16'h0392; // 0x11b2
	13'h08da: q3 = 16'hfc79; // 0x11b4
	13'h08db: q3 = 16'h8b01; // 0x11b6
	13'h08dc: q3 = 16'h0445; // 0x11b8
	13'h08dd: q3 = 16'h0400; // 0x11ba
	13'h08de: q3 = 16'h8704; // 0x11bc
	13'h08df: q3 = 16'h088b; // 0x11be
	13'h08e0: q3 = 16'h0400; // 0x11c0
	13'h08e1: q3 = 16'h8a04; // 0x11c2
	13'h08e2: q3 = 16'h0400; // 0x11c4
	13'h08e3: q3 = 16'h0a01; // 0x11c6
	13'h08e4: q3 = 16'h8e04; // 0x11c8
	13'h08e5: q3 = 16'h0000; // 0x11ca
	13'h08e6: q3 = 16'hfb46; // 0x11cc
	13'h08e7: q3 = 16'h0800; // 0x11ce
	13'h08e8: q3 = 16'h0601; // 0x11d0
	13'h08e9: q3 = 16'h0000; // 0x11d2
	13'h08ea: q3 = 16'h0000; // 0x11d4
	13'h08eb: q3 = 16'h0f00; // 0x11d6
	13'h08ec: q3 = 16'h0100; // 0x11d8
	13'h08ed: q3 = 16'h8705; // 0x11da
	13'h08ee: q3 = 16'h0199; // 0x11dc
	13'h08ef: q3 = 16'h0666; // 0x11de
	13'h08f0: q3 = 16'h0400; // 0x11e0
	13'h08f1: q3 = 16'h0701; // 0x11e2
	13'h08f2: q3 = 16'h01b1; // 0x11e4
	13'h08f3: q3 = 16'h8a04; // 0x11e6
	13'h08f4: q3 = 16'h0400; // 0x11e8
	13'h08f5: q3 = 16'h8707; // 0x11ea
	13'h08f6: q3 = 16'h0199; // 0x11ec
	13'h08f7: q3 = 16'h0222; // 0x11ee
	13'h08f8: q3 = 16'h0514; // 0x11f0
	13'h08f9: q3 = 16'h0400; // 0x11f2
	13'h08fa: q3 = 16'h0701; // 0x11f4
	13'h08fb: q3 = 16'h01b1; // 0x11f6
	13'h08fc: q3 = 16'h8a04; // 0x11f8
	13'h08fd: q3 = 16'h0400; // 0x11fa
	13'h08fe: q3 = 16'h0705; // 0x11fc
	13'h08ff: q3 = 16'h0199; // 0x11fe
	13'h0900: q3 = 16'h088b; // 0x1200
	13'h0901: q3 = 16'h8a02; // 0x1202
	13'h0902: q3 = 16'h0400; // 0x1204
	13'h0903: q3 = 16'h0701; // 0x1206
	13'h0904: q3 = 16'h01b1; // 0x1208
	13'h0905: q3 = 16'h8a04; // 0x120a
	13'h0906: q3 = 16'h0400; // 0x120c
	13'h0907: q3 = 16'h8707; // 0x120e
	13'h0908: q3 = 16'h0199; // 0x1210
	13'h0909: q3 = 16'h0222; // 0x1212
	13'h090a: q3 = 16'h0514; // 0x1214
	13'h090b: q3 = 16'h0400; // 0x1216
	13'h090c: q3 = 16'h0701; // 0x1218
	13'h090d: q3 = 16'h01b1; // 0x121a
	13'h090e: q3 = 16'h8a04; // 0x121c
	13'h090f: q3 = 16'h0400; // 0x121e
	13'h0910: q3 = 16'h0705; // 0x1220
	13'h0911: q3 = 16'h0199; // 0x1222
	13'h0912: q3 = 16'h0666; // 0x1224
	13'h0913: q3 = 16'h8a02; // 0x1226
	13'h0914: q3 = 16'h0400; // 0x1228
	13'h0915: q3 = 16'h0701; // 0x122a
	13'h0916: q3 = 16'h01b1; // 0x122c
	13'h0917: q3 = 16'h8a04; // 0x122e
	13'h0918: q3 = 16'h0400; // 0x1230
	13'h0919: q3 = 16'h8707; // 0x1232
	13'h091a: q3 = 16'h0199; // 0x1234
	13'h091b: q3 = 16'h0222; // 0x1236
	13'h091c: q3 = 16'h0514; // 0x1238
	13'h091d: q3 = 16'h0400; // 0x123a
	13'h091e: q3 = 16'h0701; // 0x123c
	13'h091f: q3 = 16'h01b1; // 0x123e
	13'h0920: q3 = 16'h8a04; // 0x1240
	13'h0921: q3 = 16'h0400; // 0x1242
	13'h0922: q3 = 16'h0705; // 0x1244
	13'h0923: q3 = 16'h0199; // 0x1246
	13'h0924: q3 = 16'h088b; // 0x1248
	13'h0925: q3 = 16'h8a02; // 0x124a
	13'h0926: q3 = 16'h0400; // 0x124c
	13'h0927: q3 = 16'h0701; // 0x124e
	13'h0928: q3 = 16'h01b1; // 0x1250
	13'h0929: q3 = 16'h8a04; // 0x1252
	13'h092a: q3 = 16'h0400; // 0x1254
	13'h092b: q3 = 16'h8707; // 0x1256
	13'h092c: q3 = 16'h0199; // 0x1258
	13'h092d: q3 = 16'h0222; // 0x125a
	13'h092e: q3 = 16'h0514; // 0x125c
	13'h092f: q3 = 16'h0400; // 0x125e
	13'h0930: q3 = 16'h0701; // 0x1260
	13'h0931: q3 = 16'h0182; // 0x1262
	13'h0932: q3 = 16'h8a04; // 0x1264
	13'h0933: q3 = 16'h0400; // 0x1266
	13'h0934: q3 = 16'h0705; // 0x1268
	13'h0935: q3 = 16'h016c; // 0x126a
	13'h0936: q3 = 16'h06c7; // 0x126c
	13'h0937: q3 = 16'h8a02; // 0x126e
	13'h0938: q3 = 16'h0400; // 0x1270
	13'h0939: q3 = 16'h8a05; // 0x1272
	13'h093a: q3 = 16'h0400; // 0x1274
	13'h093b: q3 = 16'h8707; // 0x1276
	13'h093c: q3 = 16'h01b1; // 0x1278
	13'h093d: q3 = 16'h0222; // 0x127a
	13'h093e: q3 = 16'h04cb; // 0x127c
	13'h093f: q3 = 16'h0400; // 0x127e
	13'h0940: q3 = 16'h8a05; // 0x1280
	13'h0941: q3 = 16'h0400; // 0x1282
	13'h0942: q3 = 16'h0705; // 0x1284
	13'h0943: q3 = 16'h01e7; // 0x1286
	13'h0944: q3 = 16'h088b; // 0x1288
	13'h0945: q3 = 16'h8a02; // 0x128a
	13'h0946: q3 = 16'h0400; // 0x128c
	13'h0947: q3 = 16'h0701; // 0x128e
	13'h0948: q3 = 16'h01b1; // 0x1290
	13'h0949: q3 = 16'h8a04; // 0x1292
	13'h094a: q3 = 16'h0400; // 0x1294
	13'h094b: q3 = 16'h0706; // 0x1296
	13'h094c: q3 = 16'h0222; // 0x1298
	13'h094d: q3 = 16'h04cb; // 0x129a
	13'h094e: q3 = 16'h8a01; // 0x129c
	13'h094f: q3 = 16'h0400; // 0x129e
	13'h0950: q3 = 16'h0701; // 0x12a0
	13'h0951: q3 = 16'h016c; // 0x12a2
	13'h0952: q3 = 16'h8a04; // 0x12a4
	13'h0953: q3 = 16'h0400; // 0x12a6
	13'h0954: q3 = 16'h0704; // 0x12a8
	13'h0955: q3 = 16'h06c7; // 0x12aa
	13'h0956: q3 = 16'h8a02; // 0x12ac
	13'h0957: q3 = 16'h0400; // 0x12ae
	13'h0958: q3 = 16'h8a04; // 0x12b0
	13'h0959: q3 = 16'h0400; // 0x12b2
	13'h095a: q3 = 16'h8706; // 0x12b4
	13'h095b: q3 = 16'h0222; // 0x12b6
	13'h095c: q3 = 16'h04cb; // 0x12b8
	13'h095d: q3 = 16'h0400; // 0x12ba
	13'h095e: q3 = 16'h8a04; // 0x12bc
	13'h095f: q3 = 16'h0400; // 0x12be
	13'h0960: q3 = 16'h0704; // 0x12c0
	13'h0961: q3 = 16'h088b; // 0x12c2
	13'h0962: q3 = 16'h8a02; // 0x12c4
	13'h0963: q3 = 16'h0400; // 0x12c6
	13'h0964: q3 = 16'h8a04; // 0x12c8
	13'h0965: q3 = 16'h0400; // 0x12ca
	13'h0966: q3 = 16'h8706; // 0x12cc
	13'h0967: q3 = 16'h0222; // 0x12ce
	13'h0968: q3 = 16'h04cb; // 0x12d0
	13'h0969: q3 = 16'h0400; // 0x12d2
	13'h096a: q3 = 16'h8a04; // 0x12d4
	13'h096b: q3 = 16'h0400; // 0x12d6
	13'h096c: q3 = 16'h0a03; // 0x12d8
	13'h096d: q3 = 16'h0100; // 0x12da
	13'h096e: q3 = 16'h870d; // 0x12dc
	13'h096f: q3 = 16'h01b1; // 0x12de
	13'h0970: q3 = 16'h0363; // 0x12e0
	13'h0971: q3 = 16'h05b3; // 0x12e2
	13'h0972: q3 = 16'h0400; // 0x12e4
	13'h0973: q3 = 16'h0701; // 0x12e6
	13'h0974: q3 = 16'h01cb; // 0x12e8
	13'h0975: q3 = 16'h8a04; // 0x12ea
	13'h0976: q3 = 16'h0400; // 0x12ec
	13'h0977: q3 = 16'h0707; // 0x12ee
	13'h0978: q3 = 16'h01b1; // 0x12f0
	13'h0979: q3 = 16'h0222; // 0x12f2
	13'h097a: q3 = 16'h0265; // 0x12f4
	13'h097b: q3 = 16'h8a08; // 0x12f6
	13'h097c: q3 = 16'h0400; // 0x12f8
	13'h097d: q3 = 16'h0701; // 0x12fa
	13'h097e: q3 = 16'h0222; // 0x12fc
	13'h097f: q3 = 16'h8a04; // 0x12fe
	13'h0980: q3 = 16'h0400; // 0x1300
	13'h0981: q3 = 16'h070d; // 0x1302
	13'h0982: q3 = 16'h0363; // 0x1304
	13'h0983: q3 = 16'h0445; // 0x1306
	13'h0984: q3 = 16'h088b; // 0x1308
	13'h0985: q3 = 16'h8a02; // 0x130a
	13'h0986: q3 = 16'h0400; // 0x130c
	13'h0987: q3 = 16'h0701; // 0x130e
	13'h0988: q3 = 16'h0333; // 0x1310
	13'h0989: q3 = 16'h8a04; // 0x1312
	13'h098a: q3 = 16'h0400; // 0x1314
	13'h098b: q3 = 16'h0707; // 0x1316
	13'h098c: q3 = 16'h0305; // 0x1318
	13'h098d: q3 = 16'h0222; // 0x131a
	13'h098e: q3 = 16'h0265; // 0x131c
	13'h098f: q3 = 16'h8a08; // 0x131e
	13'h0990: q3 = 16'h0400; // 0x1320
	13'h0991: q3 = 16'h0701; // 0x1322
	13'h0992: q3 = 16'h02d9; // 0x1324
	13'h0993: q3 = 16'h8a04; // 0x1326
	13'h0994: q3 = 16'h0400; // 0x1328
	13'h0995: q3 = 16'h070d; // 0x132a
	13'h0996: q3 = 16'h00d8; // 0x132c
	13'h0997: q3 = 16'h0363; // 0x132e
	13'h0998: q3 = 16'h05b3; // 0x1330
	13'h0999: q3 = 16'h8a02; // 0x1332
	13'h099a: q3 = 16'h0400; // 0x1334
	13'h099b: q3 = 16'h0701; // 0x1336
	13'h099c: q3 = 16'h00e5; // 0x1338
	13'h099d: q3 = 16'h8a04; // 0x133a
	13'h099e: q3 = 16'h0400; // 0x133c
	13'h099f: q3 = 16'h0707; // 0x133e
	13'h09a0: q3 = 16'h00f3; // 0x1340
	13'h09a1: q3 = 16'h0222; // 0x1342
	13'h09a2: q3 = 16'h0265; // 0x1344
	13'h09a3: q3 = 16'h8a08; // 0x1346
	13'h09a4: q3 = 16'h0400; // 0x1348
	13'h09a5: q3 = 16'h0701; // 0x134a
	13'h09a6: q3 = 16'h0111; // 0x134c
	13'h09a7: q3 = 16'h8a04; // 0x134e
	13'h09a8: q3 = 16'h0400; // 0x1350
	13'h09a9: q3 = 16'h070c; // 0x1352
	13'h09aa: q3 = 16'h0445; // 0x1354
	13'h09ab: q3 = 16'h088b; // 0x1356
	13'h09ac: q3 = 16'h8a02; // 0x1358
	13'h09ad: q3 = 16'h0400; // 0x135a
	13'h09ae: q3 = 16'h8a04; // 0x135c
	13'h09af: q3 = 16'h0400; // 0x135e
	13'h09b0: q3 = 16'h0705; // 0x1360
	13'h09b1: q3 = 16'h0222; // 0x1362
	13'h09b2: q3 = 16'h0265; // 0x1364
	13'h09b3: q3 = 16'h8a08; // 0x1366
	13'h09b4: q3 = 16'h0400; // 0x1368
	13'h09b5: q3 = 16'h8a04; // 0x136a
	13'h09b6: q3 = 16'h0400; // 0x136c
	13'h09b7: q3 = 16'h870d; // 0x136e
	13'h09b8: q3 = 16'h0199; // 0x1370
	13'h09b9: q3 = 16'h0333; // 0x1372
	13'h09ba: q3 = 16'h0666; // 0x1374
	13'h09bb: q3 = 16'h0400; // 0x1376
	13'h09bc: q3 = 16'h0701; // 0x1378
	13'h09bd: q3 = 16'h01b1; // 0x137a
	13'h09be: q3 = 16'h8a04; // 0x137c
	13'h09bf: q3 = 16'h0400; // 0x137e
	13'h09c0: q3 = 16'h0707; // 0x1380
	13'h09c1: q3 = 16'h0199; // 0x1382
	13'h09c2: q3 = 16'h0222; // 0x1384
	13'h09c3: q3 = 16'h028a; // 0x1386
	13'h09c4: q3 = 16'h8a08; // 0x1388
	13'h09c5: q3 = 16'h0400; // 0x138a
	13'h09c6: q3 = 16'h0701; // 0x138c
	13'h09c7: q3 = 16'h0222; // 0x138e
	13'h09c8: q3 = 16'h8a04; // 0x1390
	13'h09c9: q3 = 16'h0400; // 0x1392
	13'h09ca: q3 = 16'h070d; // 0x1394
	13'h09cb: q3 = 16'h0333; // 0x1396
	13'h09cc: q3 = 16'h0445; // 0x1398
	13'h09cd: q3 = 16'h088b; // 0x139a
	13'h09ce: q3 = 16'h8a02; // 0x139c
	13'h09cf: q3 = 16'h0400; // 0x139e
	13'h09d0: q3 = 16'h0701; // 0x13a0
	13'h09d1: q3 = 16'h02d9; // 0x13a2
	13'h09d2: q3 = 16'h8a04; // 0x13a4
	13'h09d3: q3 = 16'h0400; // 0x13a6
	13'h09d4: q3 = 16'h0707; // 0x13a8
	13'h09d5: q3 = 16'h02b0; // 0x13aa
	13'h09d6: q3 = 16'h0222; // 0x13ac
	13'h09d7: q3 = 16'h028a; // 0x13ae
	13'h09d8: q3 = 16'h8a08; // 0x13b0
	13'h09d9: q3 = 16'h0400; // 0x13b2
	13'h09da: q3 = 16'h0701; // 0x13b4
	13'h09db: q3 = 16'h028a; // 0x13b6
	13'h09dc: q3 = 16'h8a04; // 0x13b8
	13'h09dd: q3 = 16'h0400; // 0x13ba
	13'h09de: q3 = 16'h070d; // 0x13bc
	13'h09df: q3 = 16'h00cc; // 0x13be
	13'h09e0: q3 = 16'h0333; // 0x13c0
	13'h09e1: q3 = 16'h0666; // 0x13c2
	13'h09e2: q3 = 16'h8a02; // 0x13c4
	13'h09e3: q3 = 16'h0400; // 0x13c6
	13'h09e4: q3 = 16'h0701; // 0x13c8
	13'h09e5: q3 = 16'h00d8; // 0x13ca
	13'h09e6: q3 = 16'h8a04; // 0x13cc
	13'h09e7: q3 = 16'h0400; // 0x13ce
	13'h09e8: q3 = 16'h0707; // 0x13d0
	13'h09e9: q3 = 16'h00cc; // 0x13d2
	13'h09ea: q3 = 16'h0222; // 0x13d4
	13'h09eb: q3 = 16'h028a; // 0x13d6
	13'h09ec: q3 = 16'h8a08; // 0x13d8
	13'h09ed: q3 = 16'h0400; // 0x13da
	13'h09ee: q3 = 16'h0701; // 0x13dc
	13'h09ef: q3 = 16'h0111; // 0x13de
	13'h09f0: q3 = 16'h8a04; // 0x13e0
	13'h09f1: q3 = 16'h0400; // 0x13e2
	13'h09f2: q3 = 16'h070d; // 0x13e4
	13'h09f3: q3 = 16'h0222; // 0x13e6
	13'h09f4: q3 = 16'h0445; // 0x13e8
	13'h09f5: q3 = 16'h088b; // 0x13ea
	13'h09f6: q3 = 16'h8a02; // 0x13ec
	13'h09f7: q3 = 16'h0400; // 0x13ee
	13'h09f8: q3 = 16'h0701; // 0x13f0
	13'h09f9: q3 = 16'h0204; // 0x13f2
	13'h09fa: q3 = 16'h8a04; // 0x13f4
	13'h09fb: q3 = 16'h0400; // 0x13f6
	13'h09fc: q3 = 16'h0707; // 0x13f8
	13'h09fd: q3 = 16'h01e7; // 0x13fa
	13'h09fe: q3 = 16'h0222; // 0x13fc
	13'h09ff: q3 = 16'h028a; // 0x13fe
	13'h0a00: q3 = 16'h8a08; // 0x1400
	13'h0a01: q3 = 16'h0400; // 0x1402
	13'h0a02: q3 = 16'h0701; // 0x1404
	13'h0a03: q3 = 16'h01b1; // 0x1406
	13'h0a04: q3 = 16'h8a04; // 0x1408
	13'h0a05: q3 = 16'h0400; // 0x140a
	13'h0a06: q3 = 16'h0a03; // 0x140c
	13'h0a07: q3 = 16'h0100; // 0x140e
	13'h0a08: q3 = 16'h870d; // 0x1410
	13'h0a09: q3 = 16'h0132; // 0x1412
	13'h0a0a: q3 = 16'h0363; // 0x1414
	13'h0a0b: q3 = 16'h05b3; // 0x1416
	13'h0a0c: q3 = 16'h0400; // 0x1418
	13'h0a0d: q3 = 16'h0701; // 0x141a
	13'h0a0e: q3 = 16'h0145; // 0x141c
	13'h0a0f: q3 = 16'h8a04; // 0x141e
	13'h0a10: q3 = 16'h0400; // 0x1420
	13'h0a11: q3 = 16'h0707; // 0x1422
	13'h0a12: q3 = 16'h016c; // 0x1424
	13'h0a13: q3 = 16'h0222; // 0x1426
	13'h0a14: q3 = 16'h0265; // 0x1428
	13'h0a15: q3 = 16'h8a08; // 0x142a
	13'h0a16: q3 = 16'h0400; // 0x142c
	13'h0a17: q3 = 16'h0701; // 0x142e
	13'h0a18: q3 = 16'h0199; // 0x1430
	13'h0a19: q3 = 16'h8a04; // 0x1432
	13'h0a1a: q3 = 16'h0400; // 0x1434
	13'h0a1b: q3 = 16'h070d; // 0x1436
	13'h0a1c: q3 = 16'h01b1; // 0x1438
	13'h0a1d: q3 = 16'h0445; // 0x143a
	13'h0a1e: q3 = 16'h088b; // 0x143c
	13'h0a1f: q3 = 16'h8a02; // 0x143e
	13'h0a20: q3 = 16'h0400; // 0x1440
	13'h0a21: q3 = 16'h0701; // 0x1442
	13'h0a22: q3 = 16'h01e7; // 0x1444
	13'h0a23: q3 = 16'h8a04; // 0x1446
	13'h0a24: q3 = 16'h0400; // 0x1448
	13'h0a25: q3 = 16'h0707; // 0x144a
	13'h0a26: q3 = 16'h0222; // 0x144c
	13'h0a27: q3 = 16'h0222; // 0x144e
	13'h0a28: q3 = 16'h0265; // 0x1450
	13'h0a29: q3 = 16'h8a08; // 0x1452
	13'h0a2a: q3 = 16'h0400; // 0x1454
	13'h0a2b: q3 = 16'h0701; // 0x1456
	13'h0a2c: q3 = 16'h0243; // 0x1458
	13'h0a2d: q3 = 16'h8a04; // 0x145a
	13'h0a2e: q3 = 16'h0400; // 0x145c
	13'h0a2f: q3 = 16'h070d; // 0x145e
	13'h0a30: q3 = 16'h0222; // 0x1460
	13'h0a31: q3 = 16'h0363; // 0x1462
	13'h0a32: q3 = 16'h05b3; // 0x1464
	13'h0a33: q3 = 16'h8a02; // 0x1466
	13'h0a34: q3 = 16'h0400; // 0x1468
	13'h0a35: q3 = 16'h0701; // 0x146a
	13'h0a36: q3 = 16'h01e7; // 0x146c
	13'h0a37: q3 = 16'h8a04; // 0x146e
	13'h0a38: q3 = 16'h0400; // 0x1470
	13'h0a39: q3 = 16'h0707; // 0x1472
	13'h0a3a: q3 = 16'h01cb; // 0x1474
	13'h0a3b: q3 = 16'h0222; // 0x1476
	13'h0a3c: q3 = 16'h0265; // 0x1478
	13'h0a3d: q3 = 16'h8a08; // 0x147a
	13'h0a3e: q3 = 16'h0400; // 0x147c
	13'h0a3f: q3 = 16'h0701; // 0x147e
	13'h0a40: q3 = 16'h01b1; // 0x1480
	13'h0a41: q3 = 16'h8a04; // 0x1482
	13'h0a42: q3 = 16'h0400; // 0x1484
	13'h0a43: q3 = 16'h070c; // 0x1486
	13'h0a44: q3 = 16'h0445; // 0x1488
	13'h0a45: q3 = 16'h088b; // 0x148a
	13'h0a46: q3 = 16'h8a02; // 0x148c
	13'h0a47: q3 = 16'h0400; // 0x148e
	13'h0a48: q3 = 16'h0701; // 0x1490
	13'h0a49: q3 = 16'h0222; // 0x1492
	13'h0a4a: q3 = 16'h8a04; // 0x1494
	13'h0a4b: q3 = 16'h0400; // 0x1496
	13'h0a4c: q3 = 16'h0707; // 0x1498
	13'h0a4d: q3 = 16'h01e7; // 0x149a
	13'h0a4e: q3 = 16'h0222; // 0x149c
	13'h0a4f: q3 = 16'h0265; // 0x149e
	13'h0a50: q3 = 16'h8a08; // 0x14a0
	13'h0a51: q3 = 16'h0400; // 0x14a2
	13'h0a52: q3 = 16'h0701; // 0x14a4
	13'h0a53: q3 = 16'h01b1; // 0x14a6
	13'h0a54: q3 = 16'h8a04; // 0x14a8
	13'h0a55: q3 = 16'h0400; // 0x14aa
	13'h0a56: q3 = 16'h0a03; // 0x14ac
	13'h0a57: q3 = 16'h0100; // 0x14ae
	13'h0a58: q3 = 16'h870f; // 0x14b0
	13'h0a59: q3 = 16'h0199; // 0x14b2
	13'h0a5a: q3 = 16'h0333; // 0x14b4
	13'h0a5b: q3 = 16'h0ccc; // 0x14b6
	13'h0a5c: q3 = 16'h1999; // 0x14b8
	13'h0a5d: q3 = 16'h0400; // 0x14ba
	13'h0a5e: q3 = 16'h8a05; // 0x14bc
	13'h0a5f: q3 = 16'h0400; // 0x14be
	13'h0a60: q3 = 16'h0701; // 0x14c0
	13'h0a61: q3 = 16'h01e7; // 0x14c2
	13'h0a62: q3 = 16'h8a0a; // 0x14c4
	13'h0a63: q3 = 16'h0400; // 0x14c6
	13'h0a64: q3 = 16'h8a01; // 0x14c8
	13'h0a65: q3 = 16'h0400; // 0x14ca
	13'h0a66: q3 = 16'h0701; // 0x14cc
	13'h0a67: q3 = 16'h0222; // 0x14ce
	13'h0a68: q3 = 16'h8f00; // 0x14d0
	13'h0a69: q3 = 16'h0400; // 0x14d2
	13'h0a6a: q3 = 16'h8701; // 0x14d4
	13'h0a6b: q3 = 16'h01e7; // 0x14d6
	13'h0a6c: q3 = 16'h0400; // 0x14d8
	13'h0a6d: q3 = 16'h8a01; // 0x14da
	13'h0a6e: q3 = 16'h0800; // 0x14dc
	13'h0a6f: q3 = 16'h070f; // 0x14de
	13'h0a70: q3 = 16'h0199; // 0x14e0
	13'h0a71: q3 = 16'h0333; // 0x14e2
	13'h0a72: q3 = 16'h0ccc; // 0x14e4
	13'h0a73: q3 = 16'h1999; // 0x14e6
	13'h0a74: q3 = 16'h8f00; // 0x14e8
	13'h0a75: q3 = 16'h0400; // 0x14ea
	13'h0a76: q3 = 16'h8a05; // 0x14ec
	13'h0a77: q3 = 16'h0400; // 0x14ee
	13'h0a78: q3 = 16'h0701; // 0x14f0
	13'h0a79: q3 = 16'h01e7; // 0x14f2
	13'h0a7a: q3 = 16'h8a0a; // 0x14f4
	13'h0a7b: q3 = 16'h0400; // 0x14f6
	13'h0a7c: q3 = 16'h8a01; // 0x14f8
	13'h0a7d: q3 = 16'h0400; // 0x14fa
	13'h0a7e: q3 = 16'h0701; // 0x14fc
	13'h0a7f: q3 = 16'h0222; // 0x14fe
	13'h0a80: q3 = 16'h8f00; // 0x1500
	13'h0a81: q3 = 16'h0400; // 0x1502
	13'h0a82: q3 = 16'h8701; // 0x1504
	13'h0a83: q3 = 16'h01e7; // 0x1506
	13'h0a84: q3 = 16'h0400; // 0x1508
	13'h0a85: q3 = 16'h8a01; // 0x150a
	13'h0a86: q3 = 16'h0800; // 0x150c
	13'h0a87: q3 = 16'h070f; // 0x150e
	13'h0a88: q3 = 16'h0199; // 0x1510
	13'h0a89: q3 = 16'h0333; // 0x1512
	13'h0a8a: q3 = 16'h0666; // 0x1514
	13'h0a8b: q3 = 16'h1999; // 0x1516
	13'h0a8c: q3 = 16'h8f00; // 0x1518
	13'h0a8d: q3 = 16'h0400; // 0x151a
	13'h0a8e: q3 = 16'h8a05; // 0x151c
	13'h0a8f: q3 = 16'h0400; // 0x151e
	13'h0a90: q3 = 16'h0705; // 0x1520
	13'h0a91: q3 = 16'h01e7; // 0x1522
	13'h0a92: q3 = 16'h088b; // 0x1524
	13'h0a93: q3 = 16'h8a0a; // 0x1526
	13'h0a94: q3 = 16'h0400; // 0x1528
	13'h0a95: q3 = 16'h8a05; // 0x152a
	13'h0a96: q3 = 16'h0400; // 0x152c
	13'h0a97: q3 = 16'h0302; // 0x152e
	13'h0a98: q3 = 16'h0000; // 0x1530
	13'h0a99: q3 = 16'hf332; // 0x1532
	13'h0a9a: q3 = 16'h0502; // 0x1534
	13'h0a9b: q3 = 16'h0000; // 0x1536
	13'h0a9c: q3 = 16'hf34a; // 0x1538
	13'h0a9d: q3 = 16'h8705; // 0x153a
	13'h0a9e: q3 = 16'h0222; // 0x153c
	13'h0a9f: q3 = 16'h079c; // 0x153e
	13'h0aa0: q3 = 16'h0400; // 0x1540
	13'h0aa1: q3 = 16'h0701; // 0x1542
	13'h0aa2: q3 = 16'h01e7; // 0x1544
	13'h0aa3: q3 = 16'h8a04; // 0x1546
	13'h0aa4: q3 = 16'h0400; // 0x1548
	13'h0aa5: q3 = 16'h0704; // 0x154a
	13'h0aa6: q3 = 16'h06c7; // 0x154c
	13'h0aa7: q3 = 16'h8a01; // 0x154e
	13'h0aa8: q3 = 16'h0400; // 0x1550
	13'h0aa9: q3 = 16'h0703; // 0x1552
	13'h0aaa: q3 = 16'h0199; // 0x1554
	13'h0aab: q3 = 16'h0199; // 0x1556
	13'h0aac: q3 = 16'h8a04; // 0x1558
	13'h0aad: q3 = 16'h0400; // 0x155a
	13'h0aae: q3 = 16'h8704; // 0x155c
	13'h0aaf: q3 = 16'h0666; // 0x155e
	13'h0ab0: q3 = 16'h0400; // 0x1560
	13'h0ab1: q3 = 16'h8a04; // 0x1562
	13'h0ab2: q3 = 16'h0400; // 0x1564
	13'h0ab3: q3 = 16'h0603; // 0x1566
	13'h0ab4: q3 = 16'h0479; // 0x1568
	13'h0ab5: q3 = 16'hfb9a; // 0x156a
	13'h0ab6: q3 = 16'h0479; // 0x156c
	13'h0ab7: q3 = 16'hfb9a; // 0x156e
	13'h0ab8: q3 = 16'h8b03; // 0x1570
	13'h0ab9: q3 = 16'h00c7; // 0x1572
	13'h0aba: q3 = 16'h0333; // 0x1574
	13'h0abb: q3 = 16'h0800; // 0x1576
	13'h0abc: q3 = 16'h070c; // 0x1578
	13'h0abd: q3 = 16'h0ccc; // 0x157a
	13'h0abe: q3 = 16'h1999; // 0x157c
	13'h0abf: q3 = 16'h8f00; // 0x157e
	13'h0ac0: q3 = 16'h0400; // 0x1580
	13'h0ac1: q3 = 16'h8a04; // 0x1582
	13'h0ac2: q3 = 16'h0400; // 0x1584
	13'h0ac3: q3 = 16'h8a0b; // 0x1586
	13'h0ac4: q3 = 16'h1800; // 0x1588
	13'h0ac5: q3 = 16'h0100; // 0x158a
	13'h0ac6: q3 = 16'h8705; // 0x158c
	13'h0ac7: q3 = 16'h0199; // 0x158e
	13'h0ac8: q3 = 16'h0666; // 0x1590
	13'h0ac9: q3 = 16'h0400; // 0x1592
	13'h0aca: q3 = 16'h0701; // 0x1594
	13'h0acb: q3 = 16'h01b1; // 0x1596
	13'h0acc: q3 = 16'h8a04; // 0x1598
	13'h0acd: q3 = 16'h0400; // 0x159a
	13'h0ace: q3 = 16'h8707; // 0x159c
	13'h0acf: q3 = 16'h0199; // 0x159e
	13'h0ad0: q3 = 16'h0222; // 0x15a0
	13'h0ad1: q3 = 16'h0514; // 0x15a2
	13'h0ad2: q3 = 16'h0400; // 0x15a4
	13'h0ad3: q3 = 16'h0701; // 0x15a6
	13'h0ad4: q3 = 16'h01b1; // 0x15a8
	13'h0ad5: q3 = 16'h8a04; // 0x15aa
	13'h0ad6: q3 = 16'h0400; // 0x15ac
	13'h0ad7: q3 = 16'h0705; // 0x15ae
	13'h0ad8: q3 = 16'h0199; // 0x15b0
	13'h0ad9: q3 = 16'h088b; // 0x15b2
	13'h0ada: q3 = 16'h8a02; // 0x15b4
	13'h0adb: q3 = 16'h0400; // 0x15b6
	13'h0adc: q3 = 16'h0701; // 0x15b8
	13'h0add: q3 = 16'h01b1; // 0x15ba
	13'h0ade: q3 = 16'h8a04; // 0x15bc
	13'h0adf: q3 = 16'h0400; // 0x15be
	13'h0ae0: q3 = 16'h8707; // 0x15c0
	13'h0ae1: q3 = 16'h0199; // 0x15c2
	13'h0ae2: q3 = 16'h0222; // 0x15c4
	13'h0ae3: q3 = 16'h0666; // 0x15c6
	13'h0ae4: q3 = 16'h0400; // 0x15c8
	13'h0ae5: q3 = 16'h0701; // 0x15ca
	13'h0ae6: q3 = 16'h01e7; // 0x15cc
	13'h0ae7: q3 = 16'h8a04; // 0x15ce
	13'h0ae8: q3 = 16'h0400; // 0x15d0
	13'h0ae9: q3 = 16'h0705; // 0x15d2
	13'h0aea: q3 = 16'h0222; // 0x15d4
	13'h0aeb: q3 = 16'h088b; // 0x15d6
	13'h0aec: q3 = 16'h8a02; // 0x15d8
	13'h0aed: q3 = 16'h0400; // 0x15da
	13'h0aee: q3 = 16'h0701; // 0x15dc
	13'h0aef: q3 = 16'h0243; // 0x15de
	13'h0af0: q3 = 16'h8a04; // 0x15e0
	13'h0af1: q3 = 16'h0400; // 0x15e2
	13'h0af2: q3 = 16'h8707; // 0x15e4
	13'h0af3: q3 = 16'h0222; // 0x15e6
	13'h0af4: q3 = 16'h0222; // 0x15e8
	13'h0af5: q3 = 16'h06c7; // 0x15ea
	13'h0af6: q3 = 16'h0400; // 0x15ec
	13'h0af7: q3 = 16'h0701; // 0x15ee
	13'h0af8: q3 = 16'h0243; // 0x15f0
	13'h0af9: q3 = 16'h8a04; // 0x15f2
	13'h0afa: q3 = 16'h0400; // 0x15f4
	13'h0afb: q3 = 16'h0705; // 0x15f6
	13'h0afc: q3 = 16'h0222; // 0x15f8
	13'h0afd: q3 = 16'h0b67; // 0x15fa
	13'h0afe: q3 = 16'h8a02; // 0x15fc
	13'h0aff: q3 = 16'h0400; // 0x15fe
	13'h0b00: q3 = 16'h0701; // 0x1600
	13'h0b01: q3 = 16'h0204; // 0x1602
	13'h0b02: q3 = 16'h8a04; // 0x1604
	13'h0b03: q3 = 16'h0400; // 0x1606
	13'h0b04: q3 = 16'h8707; // 0x1608
	13'h0b05: q3 = 16'h01e7; // 0x160a
	13'h0b06: q3 = 16'h0222; // 0x160c
	13'h0b07: q3 = 16'h088b; // 0x160e
	13'h0b08: q3 = 16'h0400; // 0x1610
	13'h0b09: q3 = 16'h0701; // 0x1612
	13'h0b0a: q3 = 16'h01b1; // 0x1614
	13'h0b0b: q3 = 16'h8a04; // 0x1616
	13'h0b0c: q3 = 16'h0400; // 0x1618
	13'h0b0d: q3 = 16'h0a03; // 0x161a
	13'h0b0e: q3 = 16'h0100; // 0x161c
	13'h0b0f: q3 = 16'h870f; // 0x161e
	13'h0b10: q3 = 16'h0111; // 0x1620
	13'h0b11: q3 = 16'h0445; // 0x1622
	13'h0b12: q3 = 16'h088b; // 0x1624
	13'h0b13: q3 = 16'h088b; // 0x1626
	13'h0b14: q3 = 16'h0c00; // 0x1628
	13'h0b15: q3 = 16'h8703; // 0x162a
	13'h0b16: q3 = 16'h0132; // 0x162c
	13'h0b17: q3 = 16'h0408; // 0x162e
	13'h0b18: q3 = 16'h0400; // 0x1630
	13'h0b19: q3 = 16'h0703; // 0x1632
	13'h0b1a: q3 = 16'h0145; // 0x1634
	13'h0b1b: q3 = 16'h03ce; // 0x1636
	13'h0b1c: q3 = 16'h8a08; // 0x1638
	13'h0b1d: q3 = 16'h0800; // 0x163a
	13'h0b1e: q3 = 16'h8707; // 0x163c
	13'h0b1f: q3 = 16'h016c; // 0x163e
	13'h0b20: q3 = 16'h0363; // 0x1640
	13'h0b21: q3 = 16'h088b; // 0x1642
	13'h0b22: q3 = 16'h0800; // 0x1644
	13'h0b23: q3 = 16'h0a07; // 0x1646
	13'h0b24: q3 = 16'h0100; // 0x1648
	13'h0b25: q3 = 16'h870d; // 0x164a
	13'h0b26: q3 = 16'h0199; // 0x164c
	13'h0b27: q3 = 16'h0333; // 0x164e
	13'h0b28: q3 = 16'h0666; // 0x1650
	13'h0b29: q3 = 16'h0400; // 0x1652
	13'h0b2a: q3 = 16'h0701; // 0x1654
	13'h0b2b: q3 = 16'h01b1; // 0x1656
	13'h0b2c: q3 = 16'h8a04; // 0x1658
	13'h0b2d: q3 = 16'h0400; // 0x165a
	13'h0b2e: q3 = 16'h0707; // 0x165c
	13'h0b2f: q3 = 16'h0199; // 0x165e
	13'h0b30: q3 = 16'h0222; // 0x1660
	13'h0b31: q3 = 16'h028a; // 0x1662
	13'h0b32: q3 = 16'h8a08; // 0x1664
	13'h0b33: q3 = 16'h0400; // 0x1666
	13'h0b34: q3 = 16'h0701; // 0x1668
	13'h0b35: q3 = 16'h01b1; // 0x166a
	13'h0b36: q3 = 16'h8a04; // 0x166c
	13'h0b37: q3 = 16'h0400; // 0x166e
	13'h0b38: q3 = 16'h070d; // 0x1670
	13'h0b39: q3 = 16'h0199; // 0x1672
	13'h0b3a: q3 = 16'h0445; // 0x1674
	13'h0b3b: q3 = 16'h088b; // 0x1676
	13'h0b3c: q3 = 16'h8a02; // 0x1678
	13'h0b3d: q3 = 16'h0400; // 0x167a
	13'h0b3e: q3 = 16'h0701; // 0x167c
	13'h0b3f: q3 = 16'h01b1; // 0x167e
	13'h0b40: q3 = 16'h8a04; // 0x1680
	13'h0b41: q3 = 16'h0400; // 0x1682
	13'h0b42: q3 = 16'h0707; // 0x1684
	13'h0b43: q3 = 16'h0199; // 0x1686
	13'h0b44: q3 = 16'h0222; // 0x1688
	13'h0b45: q3 = 16'h028a; // 0x168a
	13'h0b46: q3 = 16'h8a08; // 0x168c
	13'h0b47: q3 = 16'h0400; // 0x168e
	13'h0b48: q3 = 16'h0701; // 0x1690
	13'h0b49: q3 = 16'h01b1; // 0x1692
	13'h0b4a: q3 = 16'h8a04; // 0x1694
	13'h0b4b: q3 = 16'h0400; // 0x1696
	13'h0b4c: q3 = 16'h070d; // 0x1698
	13'h0b4d: q3 = 16'h0199; // 0x169a
	13'h0b4e: q3 = 16'h0333; // 0x169c
	13'h0b4f: q3 = 16'h0666; // 0x169e
	13'h0b50: q3 = 16'h8a02; // 0x16a0
	13'h0b51: q3 = 16'h0400; // 0x16a2
	13'h0b52: q3 = 16'h0701; // 0x16a4
	13'h0b53: q3 = 16'h01b1; // 0x16a6
	13'h0b54: q3 = 16'h8a04; // 0x16a8
	13'h0b55: q3 = 16'h0400; // 0x16aa
	13'h0b56: q3 = 16'h0707; // 0x16ac
	13'h0b57: q3 = 16'h0199; // 0x16ae
	13'h0b58: q3 = 16'h0222; // 0x16b0
	13'h0b59: q3 = 16'h028a; // 0x16b2
	13'h0b5a: q3 = 16'h8a08; // 0x16b4
	13'h0b5b: q3 = 16'h0400; // 0x16b6
	13'h0b5c: q3 = 16'h0701; // 0x16b8
	13'h0b5d: q3 = 16'h01b1; // 0x16ba
	13'h0b5e: q3 = 16'h8a04; // 0x16bc
	13'h0b5f: q3 = 16'h0400; // 0x16be
	13'h0b60: q3 = 16'h070d; // 0x16c0
	13'h0b61: q3 = 16'h0199; // 0x16c2
	13'h0b62: q3 = 16'h0445; // 0x16c4
	13'h0b63: q3 = 16'h088b; // 0x16c6
	13'h0b64: q3 = 16'h8a02; // 0x16c8
	13'h0b65: q3 = 16'h0400; // 0x16ca
	13'h0b66: q3 = 16'h0701; // 0x16cc
	13'h0b67: q3 = 16'h01b1; // 0x16ce
	13'h0b68: q3 = 16'h8a04; // 0x16d0
	13'h0b69: q3 = 16'h0400; // 0x16d2
	13'h0b6a: q3 = 16'h0707; // 0x16d4
	13'h0b6b: q3 = 16'h0199; // 0x16d6
	13'h0b6c: q3 = 16'h0222; // 0x16d8
	13'h0b6d: q3 = 16'h028a; // 0x16da
	13'h0b6e: q3 = 16'h8a08; // 0x16dc
	13'h0b6f: q3 = 16'h0400; // 0x16de
	13'h0b70: q3 = 16'h0701; // 0x16e0
	13'h0b71: q3 = 16'h0182; // 0x16e2
	13'h0b72: q3 = 16'h8a04; // 0x16e4
	13'h0b73: q3 = 16'h0400; // 0x16e6
	13'h0b74: q3 = 16'h070d; // 0x16e8
	13'h0b75: q3 = 16'h016c; // 0x16ea
	13'h0b76: q3 = 16'h0363; // 0x16ec
	13'h0b77: q3 = 16'h05b3; // 0x16ee
	13'h0b78: q3 = 16'h8a02; // 0x16f0
	13'h0b79: q3 = 16'h0400; // 0x16f2
	13'h0b7a: q3 = 16'h8a05; // 0x16f4
	13'h0b7b: q3 = 16'h0400; // 0x16f6
	13'h0b7c: q3 = 16'h0707; // 0x16f8
	13'h0b7d: q3 = 16'h01b1; // 0x16fa
	13'h0b7e: q3 = 16'h0222; // 0x16fc
	13'h0b7f: q3 = 16'h0265; // 0x16fe
	13'h0b80: q3 = 16'h8a08; // 0x1700
	13'h0b81: q3 = 16'h0400; // 0x1702
	13'h0b82: q3 = 16'h8a05; // 0x1704
	13'h0b83: q3 = 16'h0400; // 0x1706
	13'h0b84: q3 = 16'h070d; // 0x1708
	13'h0b85: q3 = 16'h01e7; // 0x170a
	13'h0b86: q3 = 16'h0445; // 0x170c
	13'h0b87: q3 = 16'h088b; // 0x170e
	13'h0b88: q3 = 16'h8a02; // 0x1710
	13'h0b89: q3 = 16'h0400; // 0x1712
	13'h0b8a: q3 = 16'h0701; // 0x1714
	13'h0b8b: q3 = 16'h01b1; // 0x1716
	13'h0b8c: q3 = 16'h8a04; // 0x1718
	13'h0b8d: q3 = 16'h0400; // 0x171a
	13'h0b8e: q3 = 16'h0706; // 0x171c
	13'h0b8f: q3 = 16'h0222; // 0x171e
	13'h0b90: q3 = 16'h0265; // 0x1720
	13'h0b91: q3 = 16'h8a09; // 0x1722
	13'h0b92: q3 = 16'h0400; // 0x1724
	13'h0b93: q3 = 16'h0701; // 0x1726
	13'h0b94: q3 = 16'h016c; // 0x1728
	13'h0b95: q3 = 16'h8a04; // 0x172a
	13'h0b96: q3 = 16'h0400; // 0x172c
	13'h0b97: q3 = 16'h070c; // 0x172e
	13'h0b98: q3 = 16'h0363; // 0x1730
	13'h0b99: q3 = 16'h05b3; // 0x1732
	13'h0b9a: q3 = 16'h8a02; // 0x1734
	13'h0b9b: q3 = 16'h0400; // 0x1736
	13'h0b9c: q3 = 16'h8a04; // 0x1738
	13'h0b9d: q3 = 16'h0400; // 0x173a
	13'h0b9e: q3 = 16'h0706; // 0x173c
	13'h0b9f: q3 = 16'h0222; // 0x173e
	13'h0ba0: q3 = 16'h0265; // 0x1740
	13'h0ba1: q3 = 16'h8a08; // 0x1742
	13'h0ba2: q3 = 16'h0400; // 0x1744
	13'h0ba3: q3 = 16'h8a04; // 0x1746
	13'h0ba4: q3 = 16'h0400; // 0x1748
	13'h0ba5: q3 = 16'h070c; // 0x174a
	13'h0ba6: q3 = 16'h0445; // 0x174c
	13'h0ba7: q3 = 16'h088b; // 0x174e
	13'h0ba8: q3 = 16'h8a02; // 0x1750
	13'h0ba9: q3 = 16'h0400; // 0x1752
	13'h0baa: q3 = 16'h8a04; // 0x1754
	13'h0bab: q3 = 16'h0400; // 0x1756
	13'h0bac: q3 = 16'h0706; // 0x1758
	13'h0bad: q3 = 16'h0222; // 0x175a
	13'h0bae: q3 = 16'h0265; // 0x175c
	13'h0baf: q3 = 16'h8a08; // 0x175e
	13'h0bb0: q3 = 16'h0400; // 0x1760
	13'h0bb1: q3 = 16'h8a04; // 0x1762
	13'h0bb2: q3 = 16'h0400; // 0x1764
	13'h0bb3: q3 = 16'h0a03; // 0x1766
	13'h0bb4: q3 = 16'h0100; // 0x1768
	13'h0bb5: q3 = 16'h8705; // 0x176a
	13'h0bb6: q3 = 16'h01b1; // 0x176c
	13'h0bb7: q3 = 16'h06c7; // 0x176e
	13'h0bb8: q3 = 16'h0400; // 0x1770
	13'h0bb9: q3 = 16'h0701; // 0x1772
	13'h0bba: q3 = 16'h01e7; // 0x1774
	13'h0bbb: q3 = 16'h8a04; // 0x1776
	13'h0bbc: q3 = 16'h0400; // 0x1778
	13'h0bbd: q3 = 16'h8707; // 0x177a
	13'h0bbe: q3 = 16'h01b1; // 0x177c
	13'h0bbf: q3 = 16'h0222; // 0x177e
	13'h0bc0: q3 = 16'h04cb; // 0x1780
	13'h0bc1: q3 = 16'h0400; // 0x1782
	13'h0bc2: q3 = 16'h0701; // 0x1784
	13'h0bc3: q3 = 16'h0199; // 0x1786
	13'h0bc4: q3 = 16'h8a04; // 0x1788
	13'h0bc5: q3 = 16'h0400; // 0x178a
	13'h0bc6: q3 = 16'h0705; // 0x178c
	13'h0bc7: q3 = 16'h016c; // 0x178e
	13'h0bc8: q3 = 16'h088b; // 0x1790
	13'h0bc9: q3 = 16'h8a02; // 0x1792
	13'h0bca: q3 = 16'h0400; // 0x1794
	13'h0bcb: q3 = 16'h0701; // 0x1796
	13'h0bcc: q3 = 16'h01b1; // 0x1798
	13'h0bcd: q3 = 16'h8a04; // 0x179a
	13'h0bce: q3 = 16'h0400; // 0x179c
	13'h0bcf: q3 = 16'h8707; // 0x179e
	13'h0bd0: q3 = 16'h01e7; // 0x17a0
	13'h0bd1: q3 = 16'h0222; // 0x17a2
	13'h0bd2: q3 = 16'h04cb; // 0x17a4
	13'h0bd3: q3 = 16'h0400; // 0x17a6
	13'h0bd4: q3 = 16'h0701; // 0x17a8
	13'h0bd5: q3 = 16'h0222; // 0x17aa
	13'h0bd6: q3 = 16'h8a04; // 0x17ac
	13'h0bd7: q3 = 16'h0400; // 0x17ae
	13'h0bd8: q3 = 16'h0705; // 0x17b0
	13'h0bd9: q3 = 16'h01b1; // 0x17b2
	13'h0bda: q3 = 16'h06c7; // 0x17b4
	13'h0bdb: q3 = 16'h8a02; // 0x17b6
	13'h0bdc: q3 = 16'h0400; // 0x17b8
	13'h0bdd: q3 = 16'h0701; // 0x17ba
	13'h0bde: q3 = 16'h0199; // 0x17bc
	13'h0bdf: q3 = 16'h8a04; // 0x17be
	13'h0be0: q3 = 16'h0400; // 0x17c0
	13'h0be1: q3 = 16'h8705; // 0x17c2
	13'h0be2: q3 = 16'h0182; // 0x17c4
	13'h0be3: q3 = 16'h079c; // 0x17c6
	13'h0be4: q3 = 16'h0400; // 0x17c8
	13'h0be5: q3 = 16'h0701; // 0x17ca
	13'h0be6: q3 = 16'h016c; // 0x17cc
	13'h0be7: q3 = 16'h8a04; // 0x17ce
	13'h0be8: q3 = 16'h0400; // 0x17d0
	13'h0be9: q3 = 16'h8704; // 0x17d2
	13'h0bea: q3 = 16'h06c7; // 0x17d4
	13'h0beb: q3 = 16'h0400; // 0x17d6
	13'h0bec: q3 = 16'h0701; // 0x17d8
	13'h0bed: q3 = 16'h01b1; // 0x17da
	13'h0bee: q3 = 16'h8a04; // 0x17dc
	13'h0bef: q3 = 16'h0400; // 0x17de
	13'h0bf0: q3 = 16'h8705; // 0x17e0
	13'h0bf1: q3 = 16'h01e7; // 0x17e2
	13'h0bf2: q3 = 16'h088b; // 0x17e4
	13'h0bf3: q3 = 16'h0400; // 0x17e6
	13'h0bf4: q3 = 16'h0701; // 0x17e8
	13'h0bf5: q3 = 16'h0222; // 0x17ea
	13'h0bf6: q3 = 16'h8a04; // 0x17ec
	13'h0bf7: q3 = 16'h0400; // 0x17ee
	13'h0bf8: q3 = 16'h8705; // 0x17f0
	13'h0bf9: q3 = 16'h0199; // 0x17f2
	13'h0bfa: q3 = 16'h0666; // 0x17f4
	13'h0bfb: q3 = 16'h0400; // 0x17f6
	13'h0bfc: q3 = 16'h0701; // 0x17f8
	13'h0bfd: q3 = 16'h01b1; // 0x17fa
	13'h0bfe: q3 = 16'h8a04; // 0x17fc
	13'h0bff: q3 = 16'h0400; // 0x17fe
	13'h0c00: q3 = 16'h8705; // 0x1800
	13'h0c01: q3 = 16'h0199; // 0x1802
	13'h0c02: q3 = 16'h06c7; // 0x1804
	13'h0c03: q3 = 16'h0400; // 0x1806
	13'h0c04: q3 = 16'h0701; // 0x1808
	13'h0c05: q3 = 16'h016c; // 0x180a
	13'h0c06: q3 = 16'h8a04; // 0x180c
	13'h0c07: q3 = 16'h0400; // 0x180e
	13'h0c08: q3 = 16'h8705; // 0x1810
	13'h0c09: q3 = 16'h0145; // 0x1812
	13'h0c0a: q3 = 16'h079c; // 0x1814
	13'h0c0b: q3 = 16'h0400; // 0x1816
	13'h0c0c: q3 = 16'h0701; // 0x1818
	13'h0c0d: q3 = 16'h0199; // 0x181a
	13'h0c0e: q3 = 16'h8a04; // 0x181c
	13'h0c0f: q3 = 16'h0400; // 0x181e
	13'h0c10: q3 = 16'h8705; // 0x1820
	13'h0c11: q3 = 16'h01e7; // 0x1822
	13'h0c12: q3 = 16'h06c7; // 0x1824
	13'h0c13: q3 = 16'h0400; // 0x1826
	13'h0c14: q3 = 16'h0701; // 0x1828
	13'h0c15: q3 = 16'h0222; // 0x182a
	13'h0c16: q3 = 16'h8a04; // 0x182c
	13'h0c17: q3 = 16'h0400; // 0x182e
	13'h0c18: q3 = 16'h8705; // 0x1830
	13'h0c19: q3 = 16'h0199; // 0x1832
	13'h0c1a: q3 = 16'h0666; // 0x1834
	13'h0c1b: q3 = 16'h0400; // 0x1836
	13'h0c1c: q3 = 16'h0701; // 0x1838
	13'h0c1d: q3 = 16'h016c; // 0x183a
	13'h0c1e: q3 = 16'h8a04; // 0x183c
	13'h0c1f: q3 = 16'h0400; // 0x183e
	13'h0c20: q3 = 16'h8705; // 0x1840
	13'h0c21: q3 = 16'h0158; // 0x1842
	13'h0c22: q3 = 16'h06c7; // 0x1844
	13'h0c23: q3 = 16'h0400; // 0x1846
	13'h0c24: q3 = 16'h0701; // 0x1848
	13'h0c25: q3 = 16'h0145; // 0x184a
	13'h0c26: q3 = 16'h8a04; // 0x184c
	13'h0c27: q3 = 16'h0400; // 0x184e
	13'h0c28: q3 = 16'h8705; // 0x1850
	13'h0c29: q3 = 16'h0199; // 0x1852
	13'h0c2a: q3 = 16'h0666; // 0x1854
	13'h0c2b: q3 = 16'h0400; // 0x1856
	13'h0c2c: q3 = 16'h0701; // 0x1858
	13'h0c2d: q3 = 16'h01b1; // 0x185a
	13'h0c2e: q3 = 16'h8a04; // 0x185c
	13'h0c2f: q3 = 16'h0400; // 0x185e
	13'h0c30: q3 = 16'h8705; // 0x1860
	13'h0c31: q3 = 16'h01e7; // 0x1862
	13'h0c32: q3 = 16'h088b; // 0x1864
	13'h0c33: q3 = 16'h0400; // 0x1866
	13'h0c34: q3 = 16'h0701; // 0x1868
	13'h0c35: q3 = 16'h0222; // 0x186a
	13'h0c36: q3 = 16'h8a04; // 0x186c
	13'h0c37: q3 = 16'h0400; // 0x186e
	13'h0c38: q3 = 16'h0a01; // 0x1870
	13'h0c39: q3 = 16'h0100; // 0x1872
	13'h0c3a: q3 = 16'h8705; // 0x1874
	13'h0c3b: q3 = 16'h01b1; // 0x1876
	13'h0c3c: q3 = 16'h06c7; // 0x1878
	13'h0c3d: q3 = 16'h0400; // 0x187a
	13'h0c3e: q3 = 16'h0701; // 0x187c
	13'h0c3f: q3 = 16'h0199; // 0x187e
	13'h0c40: q3 = 16'h8a04; // 0x1880
	13'h0c41: q3 = 16'h0400; // 0x1882
	13'h0c42: q3 = 16'h8707; // 0x1884
	13'h0c43: q3 = 16'h016c; // 0x1886
	13'h0c44: q3 = 16'h0222; // 0x1888
	13'h0c45: q3 = 16'h04cb; // 0x188a
	13'h0c46: q3 = 16'h0400; // 0x188c
	13'h0c47: q3 = 16'h0701; // 0x188e
	13'h0c48: q3 = 16'h0199; // 0x1890
	13'h0c49: q3 = 16'h8a04; // 0x1892
	13'h0c4a: q3 = 16'h0400; // 0x1894
	13'h0c4b: q3 = 16'h0705; // 0x1896
	13'h0c4c: q3 = 16'h01b1; // 0x1898
	13'h0c4d: q3 = 16'h088b; // 0x189a
	13'h0c4e: q3 = 16'h8a02; // 0x189c
	13'h0c4f: q3 = 16'h0400; // 0x189e
	13'h0c50: q3 = 16'h0701; // 0x18a0
	13'h0c51: q3 = 16'h01cb; // 0x18a2
	13'h0c52: q3 = 16'h8a04; // 0x18a4
	13'h0c53: q3 = 16'h0400; // 0x18a6
	13'h0c54: q3 = 16'h8707; // 0x18a8
	13'h0c55: q3 = 16'h01b1; // 0x18aa
	13'h0c56: q3 = 16'h0222; // 0x18ac
	13'h0c57: q3 = 16'h04cb; // 0x18ae
	13'h0c58: q3 = 16'h0400; // 0x18b0
	13'h0c59: q3 = 16'h0701; // 0x18b2
	13'h0c5a: q3 = 16'h01cb; // 0x18b4
	13'h0c5b: q3 = 16'h8a04; // 0x18b6
	13'h0c5c: q3 = 16'h0400; // 0x18b8
	13'h0c5d: q3 = 16'h0705; // 0x18ba
	13'h0c5e: q3 = 16'h01b1; // 0x18bc
	13'h0c5f: q3 = 16'h06c7; // 0x18be
	13'h0c60: q3 = 16'h8a02; // 0x18c0
	13'h0c61: q3 = 16'h0400; // 0x18c2
	13'h0c62: q3 = 16'h0701; // 0x18c4
	13'h0c63: q3 = 16'h0199; // 0x18c6
	13'h0c64: q3 = 16'h8a04; // 0x18c8
	13'h0c65: q3 = 16'h0400; // 0x18ca
	13'h0c66: q3 = 16'h8707; // 0x18cc
	13'h0c67: q3 = 16'h0182; // 0x18ce
	13'h0c68: q3 = 16'h0222; // 0x18d0
	13'h0c69: q3 = 16'h04cb; // 0x18d2
	13'h0c6a: q3 = 16'h0400; // 0x18d4
	13'h0c6b: q3 = 16'h0701; // 0x18d6
	13'h0c6c: q3 = 16'h016c; // 0x18d8
	13'h0c6d: q3 = 16'h8a04; // 0x18da
	13'h0c6e: q3 = 16'h0400; // 0x18dc
	13'h0c6f: q3 = 16'h0704; // 0x18de
	13'h0c70: q3 = 16'h088b; // 0x18e0
	13'h0c71: q3 = 16'h8a02; // 0x18e2
	13'h0c72: q3 = 16'h0400; // 0x18e4
	13'h0c73: q3 = 16'h0701; // 0x18e6
	13'h0c74: q3 = 16'h0132; // 0x18e8
	13'h0c75: q3 = 16'h8a04; // 0x18ea
	13'h0c76: q3 = 16'h0400; // 0x18ec
	13'h0c77: q3 = 16'h8707; // 0x18ee
	13'h0c78: q3 = 16'h0145; // 0x18f0
	13'h0c79: q3 = 16'h0222; // 0x18f2
	13'h0c7a: q3 = 16'h04cb; // 0x18f4
	13'h0c7b: q3 = 16'h0400; // 0x18f6
	13'h0c7c: q3 = 16'h0701; // 0x18f8
	13'h0c7d: q3 = 16'h016c; // 0x18fa
	13'h0c7e: q3 = 16'h8a04; // 0x18fc
	13'h0c7f: q3 = 16'h0400; // 0x18fe
	13'h0c80: q3 = 16'h0a03; // 0x1900
	13'h0c81: q3 = 16'h0100; // 0x1902
	13'h0c82: q3 = 16'h8705; // 0x1904
	13'h0c83: q3 = 16'h0199; // 0x1906
	13'h0c84: q3 = 16'h0514; // 0x1908
	13'h0c85: q3 = 16'h0400; // 0x190a
	13'h0c86: q3 = 16'h8a05; // 0x190c
	13'h0c87: q3 = 16'h0400; // 0x190e
	13'h0c88: q3 = 16'h8707; // 0x1910
	13'h0c89: q3 = 16'h01e7; // 0x1912
	13'h0c8a: q3 = 16'h0222; // 0x1914
	13'h0c8b: q3 = 16'h088b; // 0x1916
	13'h0c8c: q3 = 16'h0400; // 0x1918
	13'h0c8d: q3 = 16'h8a05; // 0x191a
	13'h0c8e: q3 = 16'h0400; // 0x191c
	13'h0c8f: q3 = 16'h0705; // 0x191e
	13'h0c90: q3 = 16'h0222; // 0x1920
	13'h0c91: q3 = 16'h079c; // 0x1922
	13'h0c92: q3 = 16'h8a02; // 0x1924
	13'h0c93: q3 = 16'h0400; // 0x1926
	13'h0c94: q3 = 16'h0701; // 0x1928
	13'h0c95: q3 = 16'h01e7; // 0x192a
	13'h0c96: q3 = 16'h8a04; // 0x192c
	13'h0c97: q3 = 16'h0400; // 0x192e
	13'h0c98: q3 = 16'h0706; // 0x1930
	13'h0c99: q3 = 16'h0222; // 0x1932
	13'h0c9a: q3 = 16'h06c7; // 0x1934
	13'h0c9b: q3 = 16'h8a01; // 0x1936
	13'h0c9c: q3 = 16'h0400; // 0x1938
	13'h0c9d: q3 = 16'h0701; // 0x193a
	13'h0c9e: q3 = 16'h0199; // 0x193c
	13'h0c9f: q3 = 16'h8a04; // 0x193e
	13'h0ca0: q3 = 16'h0400; // 0x1940
	13'h0ca1: q3 = 16'h8706; // 0x1942
	13'h0ca2: q3 = 16'h0333; // 0x1944
	13'h0ca3: q3 = 16'h0666; // 0x1946
	13'h0ca4: q3 = 16'h0800; // 0x1948
	13'h0ca5: q3 = 16'h8a04; // 0x194a
	13'h0ca6: q3 = 16'h0400; // 0x194c
	13'h0ca7: q3 = 16'h0601; // 0x194e
	13'h0ca8: q3 = 16'h05fb; // 0x1950
	13'h0ca9: q3 = 16'hfa27; // 0x1952
	13'h0caa: q3 = 16'h8b01; // 0x1954
	13'h0cab: q3 = 16'h0333; // 0x1956
	13'h0cac: q3 = 16'h0400; // 0x1958
	13'h0cad: q3 = 16'h0704; // 0x195a
	13'h0cae: q3 = 16'h0666; // 0x195c
	13'h0caf: q3 = 16'h8a02; // 0x195e
	13'h0cb0: q3 = 16'h0800; // 0x1960
	13'h0cb1: q3 = 16'h8a05; // 0x1962
	13'h0cb2: q3 = 16'h0800; // 0x1964
	13'h0cb3: q3 = 16'h0601; // 0x1966
	13'h0cb4: q3 = 16'h0000; // 0x1968
	13'h0cb5: q3 = 16'h0000; // 0x196a
	13'h0cb6: q3 = 16'h0100; // 0x196c
	13'h0cb7: q3 = 16'h870d; // 0x196e
	13'h0cb8: q3 = 16'h0158; // 0x1970
	13'h0cb9: q3 = 16'h0333; // 0x1972
	13'h0cba: q3 = 16'h0a28; // 0x1974
	13'h0cbb: q3 = 16'h0200; // 0x1976
	13'h0cbc: q3 = 16'h0601; // 0x1978
	13'h0cbd: q3 = 16'h0392; // 0x197a
	13'h0cbe: q3 = 16'hfc79; // 0x197c
	13'h0cbf: q3 = 16'h8b01; // 0x197e
	13'h0cc0: q3 = 16'h0145; // 0x1980
	13'h0cc1: q3 = 16'h0200; // 0x1982
	13'h0cc2: q3 = 16'h8a04; // 0x1984
	13'h0cc3: q3 = 16'h0400; // 0x1986
	13'h0cc4: q3 = 16'h0704; // 0x1988
	13'h0cc5: q3 = 16'h028a; // 0x198a
	13'h0cc6: q3 = 16'h8a08; // 0x198c
	13'h0cc7: q3 = 16'h0400; // 0x198e
	13'h0cc8: q3 = 16'h8a04; // 0x1990
	13'h0cc9: q3 = 16'h0400; // 0x1992
	13'h0cca: q3 = 16'h0601; // 0x1994
	13'h0ccb: q3 = 16'h0000; // 0x1996
	13'h0ccc: q3 = 16'h0000; // 0x1998
	13'h0ccd: q3 = 16'h870d; // 0x199a
	13'h0cce: q3 = 16'h01b1; // 0x199c
	13'h0ccf: q3 = 16'h0445; // 0x199e
	13'h0cd0: q3 = 16'h088b; // 0x19a0
	13'h0cd1: q3 = 16'h0200; // 0x19a2
	13'h0cd2: q3 = 16'h0601; // 0x19a4
	13'h0cd3: q3 = 16'h0392; // 0x19a6
	13'h0cd4: q3 = 16'hfc79; // 0x19a8
	13'h0cd5: q3 = 16'h8b01; // 0x19aa
	13'h0cd6: q3 = 16'h0199; // 0x19ac
	13'h0cd7: q3 = 16'h0200; // 0x19ae
	13'h0cd8: q3 = 16'h8a04; // 0x19b0
	13'h0cd9: q3 = 16'h0400; // 0x19b2
	13'h0cda: q3 = 16'h0704; // 0x19b4
	13'h0cdb: q3 = 16'h0333; // 0x19b6
	13'h0cdc: q3 = 16'h8a08; // 0x19b8
	13'h0cdd: q3 = 16'h0400; // 0x19ba
	13'h0cde: q3 = 16'h8a04; // 0x19bc
	13'h0cdf: q3 = 16'h0400; // 0x19be
	13'h0ce0: q3 = 16'h0601; // 0x19c0
	13'h0ce1: q3 = 16'h0000; // 0x19c2
	13'h0ce2: q3 = 16'h0000; // 0x19c4
	13'h0ce3: q3 = 16'h870d; // 0x19c6
	13'h0ce4: q3 = 16'h0243; // 0x19c8
	13'h0ce5: q3 = 16'h0514; // 0x19ca
	13'h0ce6: q3 = 16'h0666; // 0x19cc
	13'h0ce7: q3 = 16'h0200; // 0x19ce
	13'h0ce8: q3 = 16'h0601; // 0x19d0
	13'h0ce9: q3 = 16'h0392; // 0x19d2
	13'h0cea: q3 = 16'hfc79; // 0x19d4
	13'h0ceb: q3 = 16'h8b01; // 0x19d6
	13'h0cec: q3 = 16'h0222; // 0x19d8
	13'h0ced: q3 = 16'h0200; // 0x19da
	13'h0cee: q3 = 16'h8a04; // 0x19dc
	13'h0cef: q3 = 16'h0400; // 0x19de
	13'h0cf0: q3 = 16'h0704; // 0x19e0
	13'h0cf1: q3 = 16'h0445; // 0x19e2
	13'h0cf2: q3 = 16'h8a08; // 0x19e4
	13'h0cf3: q3 = 16'h0400; // 0x19e6
	13'h0cf4: q3 = 16'h8a04; // 0x19e8
	13'h0cf5: q3 = 16'h0400; // 0x19ea
	13'h0cf6: q3 = 16'h0601; // 0x19ec
	13'h0cf7: q3 = 16'h0000; // 0x19ee
	13'h0cf8: q3 = 16'h0000; // 0x19f0
	13'h0cf9: q3 = 16'h870d; // 0x19f2
	13'h0cfa: q3 = 16'h02b0; // 0x19f4
	13'h0cfb: q3 = 16'h0666; // 0x19f6
	13'h0cfc: q3 = 16'h088b; // 0x19f8
	13'h0cfd: q3 = 16'h0200; // 0x19fa
	13'h0cfe: q3 = 16'h0601; // 0x19fc
	13'h0cff: q3 = 16'h0392; // 0x19fe
	13'h0d00: q3 = 16'hfc79; // 0x1a00
	13'h0d01: q3 = 16'h8b01; // 0x1a02
	13'h0d02: q3 = 16'h028a; // 0x1a04
	13'h0d03: q3 = 16'h0200; // 0x1a06
	13'h0d04: q3 = 16'h8a04; // 0x1a08
	13'h0d05: q3 = 16'h0400; // 0x1a0a
	13'h0d06: q3 = 16'h0704; // 0x1a0c
	13'h0d07: q3 = 16'h0514; // 0x1a0e
	13'h0d08: q3 = 16'h8a08; // 0x1a10
	13'h0d09: q3 = 16'h0400; // 0x1a12
	13'h0d0a: q3 = 16'h8a04; // 0x1a14
	13'h0d0b: q3 = 16'h0400; // 0x1a16
	13'h0d0c: q3 = 16'h0601; // 0x1a18
	13'h0d0d: q3 = 16'h0000; // 0x1a1a
	13'h0d0e: q3 = 16'h0000; // 0x1a1c
	13'h0d0f: q3 = 16'h870d; // 0x1a1e
	13'h0d10: q3 = 16'h0363; // 0x1a20
	13'h0d11: q3 = 16'h04cb; // 0x1a22
	13'h0d12: q3 = 16'h0b67; // 0x1a24
	13'h0d13: q3 = 16'h0400; // 0x1a26
	13'h0d14: q3 = 16'h0601; // 0x1a28
	13'h0d15: q3 = 16'h0c1b; // 0x1a2a
	13'h0d16: q3 = 16'hf470; // 0x1a2c
	13'h0d17: q3 = 16'h0b01; // 0x1a2e
	13'h0d18: q3 = 16'h0333; // 0x1a30
	13'h0d19: q3 = 16'h8a04; // 0x1a32
	13'h0d1a: q3 = 16'h0400; // 0x1a34
	13'h0d1b: q3 = 16'h0704; // 0x1a36
	13'h0d1c: q3 = 16'h0445; // 0x1a38
	13'h0d1d: q3 = 16'h0b01; // 0x1a3a
	13'h0d1e: q3 = 16'h02d9; // 0x1a3c
	13'h0d1f: q3 = 16'h8a08; // 0x1a3e
	13'h0d20: q3 = 16'h0400; // 0x1a40
	13'h0d21: q3 = 16'h0b01; // 0x1a42
	13'h0d22: q3 = 16'h028a; // 0x1a44
	13'h0d23: q3 = 16'h8a04; // 0x1a46
	13'h0d24: q3 = 16'h0400; // 0x1a48
	13'h0d25: q3 = 16'h070c; // 0x1a4a
	13'h0d26: q3 = 16'h06c7; // 0x1a4c
	13'h0d27: q3 = 16'h088b; // 0x1a4e
	13'h0d28: q3 = 16'h8b01; // 0x1a50
	13'h0d29: q3 = 16'h0265; // 0x1a52
	13'h0d2a: q3 = 16'h0400; // 0x1a54
	13'h0d2b: q3 = 16'h0b01; // 0x1a56
	13'h0d2c: q3 = 16'h028a; // 0x1a58
	13'h0d2d: q3 = 16'h8a04; // 0x1a5a
	13'h0d2e: q3 = 16'h0400; // 0x1a5c
	13'h0d2f: q3 = 16'h0704; // 0x1a5e
	13'h0d30: q3 = 16'h04cb; // 0x1a60
	13'h0d31: q3 = 16'h0b01; // 0x1a62
	13'h0d32: q3 = 16'h0265; // 0x1a64
	13'h0d33: q3 = 16'h8a08; // 0x1a66
	13'h0d34: q3 = 16'h0400; // 0x1a68
	13'h0d35: q3 = 16'h0b01; // 0x1a6a
	13'h0d36: q3 = 16'h028a; // 0x1a6c
	13'h0d37: q3 = 16'h8a04; // 0x1a6e
	13'h0d38: q3 = 16'h0400; // 0x1a70
	13'h0d39: q3 = 16'h070c; // 0x1a72
	13'h0d3a: q3 = 16'h05b3; // 0x1a74
	13'h0d3b: q3 = 16'h06c7; // 0x1a76
	13'h0d3c: q3 = 16'h8b01; // 0x1a78
	13'h0d3d: q3 = 16'h0265; // 0x1a7a
	13'h0d3e: q3 = 16'h0400; // 0x1a7c
	13'h0d3f: q3 = 16'h8a04; // 0x1a7e
	13'h0d40: q3 = 16'h0400; // 0x1a80
	13'h0d41: q3 = 16'h0704; // 0x1a82
	13'h0d42: q3 = 16'h04cb; // 0x1a84
	13'h0d43: q3 = 16'h8a08; // 0x1a86
	13'h0d44: q3 = 16'h0400; // 0x1a88
	13'h0d45: q3 = 16'h8a04; // 0x1a8a
	13'h0d46: q3 = 16'h0400; // 0x1a8c
	13'h0d47: q3 = 16'h870c; // 0x1a8e
	13'h0d48: q3 = 16'h088b; // 0x1a90
	13'h0d49: q3 = 16'h088b; // 0x1a92
	13'h0d4a: q3 = 16'h0400; // 0x1a94
	13'h0d4b: q3 = 16'h8a04; // 0x1a96
	13'h0d4c: q3 = 16'h0400; // 0x1a98
	13'h0d4d: q3 = 16'h0704; // 0x1a9a
	13'h0d4e: q3 = 16'h04cb; // 0x1a9c
	13'h0d4f: q3 = 16'h8a08; // 0x1a9e
	13'h0d50: q3 = 16'h0400; // 0x1aa0
	13'h0d51: q3 = 16'h8a04; // 0x1aa2
	13'h0d52: q3 = 16'h0400; // 0x1aa4
	13'h0d53: q3 = 16'h0601; // 0x1aa6
	13'h0d54: q3 = 16'h0000; // 0x1aa8
	13'h0d55: q3 = 16'h0000; // 0x1aaa
	13'h0d56: q3 = 16'h870d; // 0x1aac
	13'h0d57: q3 = 16'h0182; // 0x1aae
	13'h0d58: q3 = 16'h0363; // 0x1ab0
	13'h0d59: q3 = 16'h0b67; // 0x1ab2
	13'h0d5a: q3 = 16'h0200; // 0x1ab4
	13'h0d5b: q3 = 16'h0601; // 0x1ab6
	13'h0d5c: q3 = 16'h0392; // 0x1ab8
	13'h0d5d: q3 = 16'hfc79; // 0x1aba
	13'h0d5e: q3 = 16'h8b01; // 0x1abc
	13'h0d5f: q3 = 16'h016c; // 0x1abe
	13'h0d60: q3 = 16'h0200; // 0x1ac0
	13'h0d61: q3 = 16'h8a04; // 0x1ac2
	13'h0d62: q3 = 16'h0400; // 0x1ac4
	13'h0d63: q3 = 16'h0704; // 0x1ac6
	13'h0d64: q3 = 16'h02d9; // 0x1ac8
	13'h0d65: q3 = 16'h8a08; // 0x1aca
	13'h0d66: q3 = 16'h0400; // 0x1acc
	13'h0d67: q3 = 16'h8a04; // 0x1ace
	13'h0d68: q3 = 16'h0400; // 0x1ad0
	13'h0d69: q3 = 16'h0601; // 0x1ad2
	13'h0d6a: q3 = 16'h0000; // 0x1ad4
	13'h0d6b: q3 = 16'h0000; // 0x1ad6
	13'h0d6c: q3 = 16'h870d; // 0x1ad8
	13'h0d6d: q3 = 16'h01cb; // 0x1ada
	13'h0d6e: q3 = 16'h0445; // 0x1adc
	13'h0d6f: q3 = 16'h088b; // 0x1ade
	13'h0d70: q3 = 16'h0200; // 0x1ae0
	13'h0d71: q3 = 16'h0601; // 0x1ae2
	13'h0d72: q3 = 16'h0392; // 0x1ae4
	13'h0d73: q3 = 16'hfc79; // 0x1ae6
	13'h0d74: q3 = 16'h8b01; // 0x1ae8
	13'h0d75: q3 = 16'h01b1; // 0x1aea
	13'h0d76: q3 = 16'h0200; // 0x1aec
	13'h0d77: q3 = 16'h8a04; // 0x1aee
	13'h0d78: q3 = 16'h0400; // 0x1af0
	13'h0d79: q3 = 16'h0704; // 0x1af2
	13'h0d7a: q3 = 16'h0363; // 0x1af4
	13'h0d7b: q3 = 16'h8a08; // 0x1af6
	13'h0d7c: q3 = 16'h0400; // 0x1af8
	13'h0d7d: q3 = 16'h8a04; // 0x1afa
	13'h0d7e: q3 = 16'h0400; // 0x1afc
	13'h0d7f: q3 = 16'h0601; // 0x1afe
	13'h0d80: q3 = 16'h0000; // 0x1b00
	13'h0d81: q3 = 16'h0000; // 0x1b02
	13'h0d82: q3 = 16'h870d; // 0x1b04
	13'h0d83: q3 = 16'h0243; // 0x1b06
	13'h0d84: q3 = 16'h05b3; // 0x1b08
	13'h0d85: q3 = 16'h06c7; // 0x1b0a
	13'h0d86: q3 = 16'h0200; // 0x1b0c
	13'h0d87: q3 = 16'h0601; // 0x1b0e
	13'h0d88: q3 = 16'h0392; // 0x1b10
	13'h0d89: q3 = 16'hfc79; // 0x1b12
	13'h0d8a: q3 = 16'h8b01; // 0x1b14
	13'h0d8b: q3 = 16'h0222; // 0x1b16
	13'h0d8c: q3 = 16'h0200; // 0x1b18
	13'h0d8d: q3 = 16'h8a04; // 0x1b1a
	13'h0d8e: q3 = 16'h0400; // 0x1b1c
	13'h0d8f: q3 = 16'h0704; // 0x1b1e
	13'h0d90: q3 = 16'h0445; // 0x1b20
	13'h0d91: q3 = 16'h8a08; // 0x1b22
	13'h0d92: q3 = 16'h0400; // 0x1b24
	13'h0d93: q3 = 16'h8a04; // 0x1b26
	13'h0d94: q3 = 16'h0400; // 0x1b28
	13'h0d95: q3 = 16'h0601; // 0x1b2a
	13'h0d96: q3 = 16'h0000; // 0x1b2c
	13'h0d97: q3 = 16'h0000; // 0x1b2e
	13'h0d98: q3 = 16'h870d; // 0x1b30
	13'h0d99: q3 = 16'h0397; // 0x1b32
	13'h0d9a: q3 = 16'h05b3; // 0x1b34
	13'h0d9b: q3 = 16'h088b; // 0x1b36
	13'h0d9c: q3 = 16'h0200; // 0x1b38
	13'h0d9d: q3 = 16'h0601; // 0x1b3a
	13'h0d9e: q3 = 16'h0392; // 0x1b3c
	13'h0d9f: q3 = 16'hfc79; // 0x1b3e
	13'h0da0: q3 = 16'h8b01; // 0x1b40
	13'h0da1: q3 = 16'h0363; // 0x1b42
	13'h0da2: q3 = 16'h0200; // 0x1b44
	13'h0da3: q3 = 16'h8a04; // 0x1b46
	13'h0da4: q3 = 16'h0400; // 0x1b48
	13'h0da5: q3 = 16'h0704; // 0x1b4a
	13'h0da6: q3 = 16'h06c7; // 0x1b4c
	13'h0da7: q3 = 16'h8a08; // 0x1b4e
	13'h0da8: q3 = 16'h0400; // 0x1b50
	13'h0da9: q3 = 16'h8a04; // 0x1b52
	13'h0daa: q3 = 16'h0400; // 0x1b54
	13'h0dab: q3 = 16'h0601; // 0x1b56
	13'h0dac: q3 = 16'h0000; // 0x1b58
	13'h0dad: q3 = 16'h0000; // 0x1b5a
	13'h0dae: q3 = 16'h870d; // 0x1b5c
	13'h0daf: q3 = 16'h0333; // 0x1b5e
	13'h0db0: q3 = 16'h0666; // 0x1b60
	13'h0db1: q3 = 16'h0ccc; // 0x1b62
	13'h0db2: q3 = 16'h0400; // 0x1b64
	13'h0db3: q3 = 16'h0601; // 0x1b66
	13'h0db4: q3 = 16'h0c1b; // 0x1b68
	13'h0db5: q3 = 16'hf470; // 0x1b6a
	13'h0db6: q3 = 16'h0b01; // 0x1b6c
	13'h0db7: q3 = 16'h0363; // 0x1b6e
	13'h0db8: q3 = 16'h8a04; // 0x1b70
	13'h0db9: q3 = 16'h0400; // 0x1b72
	13'h0dba: q3 = 16'h0704; // 0x1b74
	13'h0dbb: q3 = 16'h0514; // 0x1b76
	13'h0dbc: q3 = 16'h0b01; // 0x1b78
	13'h0dbd: q3 = 16'h0333; // 0x1b7a
	13'h0dbe: q3 = 16'h8a08; // 0x1b7c
	13'h0dbf: q3 = 16'h0400; // 0x1b7e
	13'h0dc0: q3 = 16'h0601; // 0x1b80
	13'h0dc1: q3 = 16'h0000; // 0x1b82
	13'h0dc2: q3 = 16'h0000; // 0x1b84
	13'h0dc3: q3 = 16'h0701; // 0x1b86
	13'h0dc4: q3 = 16'h0445; // 0x1b88
	13'h0dc5: q3 = 16'h8a04; // 0x1b8a
	13'h0dc6: q3 = 16'h0400; // 0x1b8c
	13'h0dc7: q3 = 16'h870d; // 0x1b8e
	13'h0dc8: q3 = 16'h028a; // 0x1b90
	13'h0dc9: q3 = 16'h0445; // 0x1b92
	13'h0dca: q3 = 16'h088b; // 0x1b94
	13'h0dcb: q3 = 16'h0400; // 0x1b96
	13'h0dcc: q3 = 16'h0601; // 0x1b98
	13'h0dcd: q3 = 16'h0c1b; // 0x1b9a
	13'h0dce: q3 = 16'hf470; // 0x1b9c
	13'h0dcf: q3 = 16'h0b01; // 0x1b9e
	13'h0dd0: q3 = 16'h02b0; // 0x1ba0
	13'h0dd1: q3 = 16'h8a04; // 0x1ba2
	13'h0dd2: q3 = 16'h0400; // 0x1ba4
	13'h0dd3: q3 = 16'h0704; // 0x1ba6
	13'h0dd4: q3 = 16'h0514; // 0x1ba8
	13'h0dd5: q3 = 16'h0b01; // 0x1baa
	13'h0dd6: q3 = 16'h028a; // 0x1bac
	13'h0dd7: q3 = 16'h8a08; // 0x1bae
	13'h0dd8: q3 = 16'h0400; // 0x1bb0
	13'h0dd9: q3 = 16'h0601; // 0x1bb2
	13'h0dda: q3 = 16'h0000; // 0x1bb4
	13'h0ddb: q3 = 16'h0000; // 0x1bb6
	13'h0ddc: q3 = 16'h0701; // 0x1bb8
	13'h0ddd: q3 = 16'h0333; // 0x1bba
	13'h0dde: q3 = 16'h8a04; // 0x1bbc
	13'h0ddf: q3 = 16'h0400; // 0x1bbe
	13'h0de0: q3 = 16'h870d; // 0x1bc0
	13'h0de1: q3 = 16'h0222; // 0x1bc2
	13'h0de2: q3 = 16'h0666; // 0x1bc4
	13'h0de3: q3 = 16'h0514; // 0x1bc6
	13'h0de4: q3 = 16'h0400; // 0x1bc8
	13'h0de5: q3 = 16'h0601; // 0x1bca
	13'h0de6: q3 = 16'h0c1b; // 0x1bcc
	13'h0de7: q3 = 16'hf470; // 0x1bce
	13'h0de8: q3 = 16'h0b01; // 0x1bd0
	13'h0de9: q3 = 16'h0243; // 0x1bd2
	13'h0dea: q3 = 16'h8a04; // 0x1bd4
	13'h0deb: q3 = 16'h0400; // 0x1bd6
	13'h0dec: q3 = 16'h0704; // 0x1bd8
	13'h0ded: q3 = 16'h0514; // 0x1bda
	13'h0dee: q3 = 16'h0b01; // 0x1bdc
	13'h0def: q3 = 16'h0222; // 0x1bde
	13'h0df0: q3 = 16'h8a08; // 0x1be0
	13'h0df1: q3 = 16'h0400; // 0x1be2
	13'h0df2: q3 = 16'h0601; // 0x1be4
	13'h0df3: q3 = 16'h0000; // 0x1be6
	13'h0df4: q3 = 16'h0000; // 0x1be8
	13'h0df5: q3 = 16'h0701; // 0x1bea
	13'h0df6: q3 = 16'h028a; // 0x1bec
	13'h0df7: q3 = 16'h8a04; // 0x1bee
	13'h0df8: q3 = 16'h0400; // 0x1bf0
	13'h0df9: q3 = 16'h870d; // 0x1bf2
	13'h0dfa: q3 = 16'h0199; // 0x1bf4
	13'h0dfb: q3 = 16'h0445; // 0x1bf6
	13'h0dfc: q3 = 16'h088b; // 0x1bf8
	13'h0dfd: q3 = 16'h0400; // 0x1bfa
	13'h0dfe: q3 = 16'h0601; // 0x1bfc
	13'h0dff: q3 = 16'h0c1b; // 0x1bfe
	13'h0e00: q3 = 16'hf470; // 0x1c00
	13'h0e01: q3 = 16'h0b01; // 0x1c02
	13'h0e02: q3 = 16'h01b1; // 0x1c04
	13'h0e03: q3 = 16'h8a04; // 0x1c06
	13'h0e04: q3 = 16'h0400; // 0x1c08
	13'h0e05: q3 = 16'h0704; // 0x1c0a
	13'h0e06: q3 = 16'h0514; // 0x1c0c
	13'h0e07: q3 = 16'h0b01; // 0x1c0e
	13'h0e08: q3 = 16'h0199; // 0x1c10
	13'h0e09: q3 = 16'h8a08; // 0x1c12
	13'h0e0a: q3 = 16'h0400; // 0x1c14
	13'h0e0b: q3 = 16'h0601; // 0x1c16
	13'h0e0c: q3 = 16'h0000; // 0x1c18
	13'h0e0d: q3 = 16'h0000; // 0x1c1a
	13'h0e0e: q3 = 16'h0701; // 0x1c1c
	13'h0e0f: q3 = 16'h0222; // 0x1c1e
	13'h0e10: q3 = 16'h8a04; // 0x1c20
	13'h0e11: q3 = 16'h0400; // 0x1c22
	13'h0e12: q3 = 16'h870d; // 0x1c24
	13'h0e13: q3 = 16'h0158; // 0x1c26
	13'h0e14: q3 = 16'h0333; // 0x1c28
	13'h0e15: q3 = 16'h0ccc; // 0x1c2a
	13'h0e16: q3 = 16'h0200; // 0x1c2c
	13'h0e17: q3 = 16'h0601; // 0x1c2e
	13'h0e18: q3 = 16'h0392; // 0x1c30
	13'h0e19: q3 = 16'hfc79; // 0x1c32
	13'h0e1a: q3 = 16'h8b01; // 0x1c34
	13'h0e1b: q3 = 16'h0145; // 0x1c36
	13'h0e1c: q3 = 16'h0200; // 0x1c38
	13'h0e1d: q3 = 16'h8a04; // 0x1c3a
	13'h0e1e: q3 = 16'h0400; // 0x1c3c
	13'h0e1f: q3 = 16'h0704; // 0x1c3e
	13'h0e20: q3 = 16'h028a; // 0x1c40
	13'h0e21: q3 = 16'h8a08; // 0x1c42
	13'h0e22: q3 = 16'h0400; // 0x1c44
	13'h0e23: q3 = 16'h8a04; // 0x1c46
	13'h0e24: q3 = 16'h0400; // 0x1c48
	13'h0e25: q3 = 16'h0601; // 0x1c4a
	13'h0e26: q3 = 16'h0000; // 0x1c4c
	13'h0e27: q3 = 16'h0000; // 0x1c4e
	13'h0e28: q3 = 16'h870d; // 0x1c50
	13'h0e29: q3 = 16'h01b1; // 0x1c52
	13'h0e2a: q3 = 16'h0445; // 0x1c54
	13'h0e2b: q3 = 16'h088b; // 0x1c56
	13'h0e2c: q3 = 16'h0200; // 0x1c58
	13'h0e2d: q3 = 16'h0601; // 0x1c5a
	13'h0e2e: q3 = 16'h0392; // 0x1c5c
	13'h0e2f: q3 = 16'hfc79; // 0x1c5e
	13'h0e30: q3 = 16'h8b01; // 0x1c60
	13'h0e31: q3 = 16'h0199; // 0x1c62
	13'h0e32: q3 = 16'h0200; // 0x1c64
	13'h0e33: q3 = 16'h8a04; // 0x1c66
	13'h0e34: q3 = 16'h0400; // 0x1c68
	13'h0e35: q3 = 16'h0704; // 0x1c6a
	13'h0e36: q3 = 16'h0333; // 0x1c6c
	13'h0e37: q3 = 16'h8a08; // 0x1c6e
	13'h0e38: q3 = 16'h0400; // 0x1c70
	13'h0e39: q3 = 16'h8a04; // 0x1c72
	13'h0e3a: q3 = 16'h0400; // 0x1c74
	13'h0e3b: q3 = 16'h0601; // 0x1c76
	13'h0e3c: q3 = 16'h0000; // 0x1c78
	13'h0e3d: q3 = 16'h0000; // 0x1c7a
	13'h0e3e: q3 = 16'h0302; // 0x1c7c
	13'h0e3f: q3 = 16'h0000; // 0x1c7e
	13'h0e40: q3 = 16'hf332; // 0x1c80
	13'h0e41: q3 = 16'h0502; // 0x1c82
	13'h0e42: q3 = 16'h0000; // 0x1c84
	13'h0e43: q3 = 16'hf34a; // 0x1c86
	13'h0e44: q3 = 16'h870f; // 0x1c88
	13'h0e45: q3 = 16'h0243; // 0x1c8a
	13'h0e46: q3 = 16'h0158; // 0x1c8c
	13'h0e47: q3 = 16'h0514; // 0x1c8e
	13'h0e48: q3 = 16'h0666; // 0x1c90
	13'h0e49: q3 = 16'h0200; // 0x1c92
	13'h0e4a: q3 = 16'h0603; // 0x1c94
	13'h0e4b: q3 = 16'h0392; // 0x1c96
	13'h0e4c: q3 = 16'hfc79; // 0x1c98
	13'h0e4d: q3 = 16'h0392; // 0x1c9a
	13'h0e4e: q3 = 16'hfc79; // 0x1c9c
	13'h0e4f: q3 = 16'h8b03; // 0x1c9e
	13'h0e50: q3 = 16'h0222; // 0x1ca0
	13'h0e51: q3 = 16'h0145; // 0x1ca2
	13'h0e52: q3 = 16'h0200; // 0x1ca4
	13'h0e53: q3 = 16'h8a04; // 0x1ca6
	13'h0e54: q3 = 16'h0400; // 0x1ca8
	13'h0e55: q3 = 16'h0704; // 0x1caa
	13'h0e56: q3 = 16'h0445; // 0x1cac
	13'h0e57: q3 = 16'h8a08; // 0x1cae
	13'h0e58: q3 = 16'h0400; // 0x1cb0
	13'h0e59: q3 = 16'h8a04; // 0x1cb2
	13'h0e5a: q3 = 16'h0400; // 0x1cb4
	13'h0e5b: q3 = 16'h0603; // 0x1cb6
	13'h0e5c: q3 = 16'h0000; // 0x1cb8
	13'h0e5d: q3 = 16'h0000; // 0x1cba
	13'h0e5e: q3 = 16'h0000; // 0x1cbc
	13'h0e5f: q3 = 16'h0000; // 0x1cbe
	13'h0e60: q3 = 16'h870f; // 0x1cc0
	13'h0e61: q3 = 16'h02b0; // 0x1cc2
	13'h0e62: q3 = 16'h01b1; // 0x1cc4
	13'h0e63: q3 = 16'h0666; // 0x1cc6
	13'h0e64: q3 = 16'h088b; // 0x1cc8
	13'h0e65: q3 = 16'h0200; // 0x1cca
	13'h0e66: q3 = 16'h0603; // 0x1ccc
	13'h0e67: q3 = 16'h0392; // 0x1cce
	13'h0e68: q3 = 16'hfc79; // 0x1cd0
	13'h0e69: q3 = 16'h0392; // 0x1cd2
	13'h0e6a: q3 = 16'hfc79; // 0x1cd4
	13'h0e6b: q3 = 16'h8b03; // 0x1cd6
	13'h0e6c: q3 = 16'h028a; // 0x1cd8
	13'h0e6d: q3 = 16'h0199; // 0x1cda
	13'h0e6e: q3 = 16'h0200; // 0x1cdc
	13'h0e6f: q3 = 16'h8a04; // 0x1cde
	13'h0e70: q3 = 16'h0400; // 0x1ce0
	13'h0e71: q3 = 16'h0704; // 0x1ce2
	13'h0e72: q3 = 16'h0514; // 0x1ce4
	13'h0e73: q3 = 16'h8a08; // 0x1ce6
	13'h0e74: q3 = 16'h0400; // 0x1ce8
	13'h0e75: q3 = 16'h8a04; // 0x1cea
	13'h0e76: q3 = 16'h0400; // 0x1cec
	13'h0e77: q3 = 16'h0603; // 0x1cee
	13'h0e78: q3 = 16'h0000; // 0x1cf0
	13'h0e79: q3 = 16'h0000; // 0x1cf2
	13'h0e7a: q3 = 16'h0000; // 0x1cf4
	13'h0e7b: q3 = 16'h0000; // 0x1cf6
	13'h0e7c: q3 = 16'h870f; // 0x1cf8
	13'h0e7d: q3 = 16'h0102; // 0x1cfa
	13'h0e7e: q3 = 16'h01b1; // 0x1cfc
	13'h0e7f: q3 = 16'h04cb; // 0x1cfe
	13'h0e80: q3 = 16'h0996; // 0x1d00
	13'h0e81: q3 = 16'h0200; // 0x1d02
	13'h0e82: q3 = 16'h0603; // 0x1d04
	13'h0e83: q3 = 16'h0392; // 0x1d06
	13'h0e84: q3 = 16'hfc79; // 0x1d08
	13'h0e85: q3 = 16'h0392; // 0x1d0a
	13'h0e86: q3 = 16'hfc79; // 0x1d0c
	13'h0e87: q3 = 16'h8b03; // 0x1d0e
	13'h0e88: q3 = 16'h00f3; // 0x1d10
	13'h0e89: q3 = 16'h0199; // 0x1d12
	13'h0e8a: q3 = 16'h0200; // 0x1d14
	13'h0e8b: q3 = 16'h8a04; // 0x1d16
	13'h0e8c: q3 = 16'h0400; // 0x1d18
	13'h0e8d: q3 = 16'h0704; // 0x1d1a
	13'h0e8e: q3 = 16'h03ce; // 0x1d1c
	13'h0e8f: q3 = 16'h8a08; // 0x1d1e
	13'h0e90: q3 = 16'h0400; // 0x1d20
	13'h0e91: q3 = 16'h8a04; // 0x1d22
	13'h0e92: q3 = 16'h0400; // 0x1d24
	13'h0e93: q3 = 16'h0603; // 0x1d26
	13'h0e94: q3 = 16'h0000; // 0x1d28
	13'h0e95: q3 = 16'h0000; // 0x1d2a
	13'h0e96: q3 = 16'h0000; // 0x1d2c
	13'h0e97: q3 = 16'h0000; // 0x1d2e
	13'h0e98: q3 = 16'h870f; // 0x1d30
	13'h0e99: q3 = 16'h0145; // 0x1d32
	13'h0e9a: q3 = 16'h0204; // 0x1d34
	13'h0e9b: q3 = 16'h0666; // 0x1d36
	13'h0e9c: q3 = 16'h079c; // 0x1d38
	13'h0e9d: q3 = 16'h0200; // 0x1d3a
	13'h0e9e: q3 = 16'h0603; // 0x1d3c
	13'h0e9f: q3 = 16'h0392; // 0x1d3e
	13'h0ea0: q3 = 16'hfc79; // 0x1d40
	13'h0ea1: q3 = 16'h0392; // 0x1d42
	13'h0ea2: q3 = 16'hfc79; // 0x1d44
	13'h0ea3: q3 = 16'h8b03; // 0x1d46
	13'h0ea4: q3 = 16'h0132; // 0x1d48
	13'h0ea5: q3 = 16'h0199; // 0x1d4a
	13'h0ea6: q3 = 16'h0200; // 0x1d4c
	13'h0ea7: q3 = 16'h8a04; // 0x1d4e
	13'h0ea8: q3 = 16'h0400; // 0x1d50
	13'h0ea9: q3 = 16'h0704; // 0x1d52
	13'h0eaa: q3 = 16'h04cb; // 0x1d54
	13'h0eab: q3 = 16'h8a08; // 0x1d56
	13'h0eac: q3 = 16'h0400; // 0x1d58
	13'h0ead: q3 = 16'h8a04; // 0x1d5a
	13'h0eae: q3 = 16'h0400; // 0x1d5c
	13'h0eaf: q3 = 16'h0603; // 0x1d5e
	13'h0eb0: q3 = 16'h0000; // 0x1d60
	13'h0eb1: q3 = 16'h0000; // 0x1d62
	13'h0eb2: q3 = 16'h0000; // 0x1d64
	13'h0eb3: q3 = 16'h0000; // 0x1d66
	13'h0eb4: q3 = 16'h870f; // 0x1d68
	13'h0eb5: q3 = 16'h01b1; // 0x1d6a
	13'h0eb6: q3 = 16'h028a; // 0x1d6c
	13'h0eb7: q3 = 16'h079c; // 0x1d6e
	13'h0eb8: q3 = 16'h03ce; // 0x1d70
	13'h0eb9: q3 = 16'h0200; // 0x1d72
	13'h0eba: q3 = 16'h0603; // 0x1d74
	13'h0ebb: q3 = 16'h0392; // 0x1d76
	13'h0ebc: q3 = 16'hfc79; // 0x1d78
	13'h0ebd: q3 = 16'h0392; // 0x1d7a
	13'h0ebe: q3 = 16'hfc79; // 0x1d7c
	13'h0ebf: q3 = 16'h8b03; // 0x1d7e
	13'h0ec0: q3 = 16'h0199; // 0x1d80
	13'h0ec1: q3 = 16'h0265; // 0x1d82
	13'h0ec2: q3 = 16'h0200; // 0x1d84
	13'h0ec3: q3 = 16'h8a04; // 0x1d86
	13'h0ec4: q3 = 16'h0400; // 0x1d88
	13'h0ec5: q3 = 16'h0704; // 0x1d8a
	13'h0ec6: q3 = 16'h0666; // 0x1d8c
	13'h0ec7: q3 = 16'h8a08; // 0x1d8e
	13'h0ec8: q3 = 16'h0400; // 0x1d90
	13'h0ec9: q3 = 16'h8a04; // 0x1d92
	13'h0eca: q3 = 16'h0400; // 0x1d94
	13'h0ecb: q3 = 16'h0603; // 0x1d96
	13'h0ecc: q3 = 16'h0000; // 0x1d98
	13'h0ecd: q3 = 16'h0000; // 0x1d9a
	13'h0ece: q3 = 16'h0000; // 0x1d9c
	13'h0ecf: q3 = 16'h0000; // 0x1d9e
	13'h0ed0: q3 = 16'h870f; // 0x1da0
	13'h0ed1: q3 = 16'h0204; // 0x1da2
	13'h0ed2: q3 = 16'h0363; // 0x1da4
	13'h0ed3: q3 = 16'h0996; // 0x1da6
	13'h0ed4: q3 = 16'h0666; // 0x1da8
	13'h0ed5: q3 = 16'h0200; // 0x1daa
	13'h0ed6: q3 = 16'h0603; // 0x1dac
	13'h0ed7: q3 = 16'h0392; // 0x1dae
	13'h0ed8: q3 = 16'hfc79; // 0x1db0
	13'h0ed9: q3 = 16'h0392; // 0x1db2
	13'h0eda: q3 = 16'hfc79; // 0x1db4
	13'h0edb: q3 = 16'h8b03; // 0x1db6
	13'h0edc: q3 = 16'h01e7; // 0x1db8
	13'h0edd: q3 = 16'h0333; // 0x1dba
	13'h0ede: q3 = 16'h0200; // 0x1dbc
	13'h0edf: q3 = 16'h8a04; // 0x1dbe
	13'h0ee0: q3 = 16'h0400; // 0x1dc0
	13'h0ee1: q3 = 16'h0704; // 0x1dc2
	13'h0ee2: q3 = 16'h079c; // 0x1dc4
	13'h0ee3: q3 = 16'h8a08; // 0x1dc6
	13'h0ee4: q3 = 16'h0400; // 0x1dc8
	13'h0ee5: q3 = 16'h8a04; // 0x1dca
	13'h0ee6: q3 = 16'h0400; // 0x1dcc
	13'h0ee7: q3 = 16'h0603; // 0x1dce
	13'h0ee8: q3 = 16'h0000; // 0x1dd0
	13'h0ee9: q3 = 16'h0000; // 0x1dd2
	13'h0eea: q3 = 16'h0000; // 0x1dd4
	13'h0eeb: q3 = 16'h0000; // 0x1dd6
	13'h0eec: q3 = 16'h870f; // 0x1dd8
	13'h0eed: q3 = 16'h0102; // 0x1dda
	13'h0eee: q3 = 16'h0204; // 0x1ddc
	13'h0eef: q3 = 16'h0810; // 0x1dde
	13'h0ef0: q3 = 16'h0666; // 0x1de0
	13'h0ef1: q3 = 16'h0400; // 0x1de2
	13'h0ef2: q3 = 16'h0701; // 0x1de4
	13'h0ef3: q3 = 16'h0158; // 0x1de6
	13'h0ef4: q3 = 16'h8a06; // 0x1de8
	13'h0ef5: q3 = 16'h0400; // 0x1dea
	13'h0ef6: q3 = 16'h8703; // 0x1dec
	13'h0ef7: q3 = 16'h0199; // 0x1dee
	13'h0ef8: q3 = 16'h02b0; // 0x1df0
	13'h0ef9: q3 = 16'h0400; // 0x1df2
	13'h0efa: q3 = 16'h0701; // 0x1df4
	13'h0efb: q3 = 16'h0204; // 0x1df6
	13'h0efc: q3 = 16'h8a02; // 0x1df8
	13'h0efd: q3 = 16'h0400; // 0x1dfa
	13'h0efe: q3 = 16'h8702; // 0x1dfc
	13'h0eff: q3 = 16'h0333; // 0x1dfe
	13'h0f00: q3 = 16'h0400; // 0x1e00
	13'h0f01: q3 = 16'h8703; // 0x1e02
	13'h0f02: q3 = 16'h0199; // 0x1e04
	13'h0f03: q3 = 16'h0204; // 0x1e06
	13'h0f04: q3 = 16'h0199; // 0x1e08
	13'h0f05: q3 = 16'h8a08; // 0x1e0a
	13'h0f06: q3 = 16'h0267; // 0x1e0c
	13'h0f07: q3 = 16'h070d; // 0x1e0e
	13'h0f08: q3 = 16'h0158; // 0x1e10
	13'h0f09: q3 = 16'h0810; // 0x1e12
	13'h0f0a: q3 = 16'h0666; // 0x1e14
	13'h0f0b: q3 = 16'h8a02; // 0x1e16
	13'h0f0c: q3 = 16'h0400; // 0x1e18
	13'h0f0d: q3 = 16'h0701; // 0x1e1a
	13'h0f0e: q3 = 16'h0102; // 0x1e1c
	13'h0f0f: q3 = 16'h8a04; // 0x1e1e
	13'h0f10: q3 = 16'h0333; // 0x1e20
	13'h0f11: q3 = 16'h8a08; // 0x1e22
	13'h0f12: q3 = 16'h00cd; // 0x1e24
	13'h0f13: q3 = 16'h870f; // 0x1e26
	13'h0f14: q3 = 16'h0111; // 0x1e28
	13'h0f15: q3 = 16'h0222; // 0x1e2a
	13'h0f16: q3 = 16'h088b; // 0x1e2c
	13'h0f17: q3 = 16'h0666; // 0x1e2e
	13'h0f18: q3 = 16'h0400; // 0x1e30
	13'h0f19: q3 = 16'h0701; // 0x1e32
	13'h0f1a: q3 = 16'h0145; // 0x1e34
	13'h0f1b: q3 = 16'h8a06; // 0x1e36
	13'h0f1c: q3 = 16'h0400; // 0x1e38
	13'h0f1d: q3 = 16'h8703; // 0x1e3a
	13'h0f1e: q3 = 16'h0199; // 0x1e3c
	13'h0f1f: q3 = 16'h028a; // 0x1e3e
	13'h0f20: q3 = 16'h0400; // 0x1e40
	13'h0f21: q3 = 16'h0701; // 0x1e42
	13'h0f22: q3 = 16'h0222; // 0x1e44
	13'h0f23: q3 = 16'h8a02; // 0x1e46
	13'h0f24: q3 = 16'h0400; // 0x1e48
	13'h0f25: q3 = 16'h8702; // 0x1e4a
	13'h0f26: q3 = 16'h0333; // 0x1e4c
	13'h0f27: q3 = 16'h0400; // 0x1e4e
	13'h0f28: q3 = 16'h8703; // 0x1e50
	13'h0f29: q3 = 16'h0199; // 0x1e52
	13'h0f2a: q3 = 16'h028a; // 0x1e54
	13'h0f2b: q3 = 16'h0199; // 0x1e56
	13'h0f2c: q3 = 16'h8a08; // 0x1e58
	13'h0f2d: q3 = 16'h0267; // 0x1e5a
	13'h0f2e: q3 = 16'h0709; // 0x1e5c
	13'h0f2f: q3 = 16'h0145; // 0x1e5e
	13'h0f30: q3 = 16'h0666; // 0x1e60
	13'h0f31: q3 = 16'h8a02; // 0x1e62
	13'h0f32: q3 = 16'h0400; // 0x1e64
	13'h0f33: q3 = 16'h8701; // 0x1e66
	13'h0f34: q3 = 16'h0132; // 0x1e68
	13'h0f35: q3 = 16'h0333; // 0x1e6a
	13'h0f36: q3 = 16'h8a08; // 0x1e6c
	13'h0f37: q3 = 16'h00cd; // 0x1e6e
	13'h0f38: q3 = 16'h870f; // 0x1e70
	13'h0f39: q3 = 16'h0111; // 0x1e72
	13'h0f3a: q3 = 16'h0445; // 0x1e74
	13'h0f3b: q3 = 16'h088b; // 0x1e76
	13'h0f3c: q3 = 16'h0445; // 0x1e78
	13'h0f3d: q3 = 16'h0600; // 0x1e7a
	13'h0f3e: q3 = 16'h8a01; // 0x1e7c
	13'h0f3f: q3 = 16'h0600; // 0x1e7e
	13'h0f40: q3 = 16'h0703; // 0x1e80
	13'h0f41: q3 = 16'h0132; // 0x1e82
	13'h0f42: q3 = 16'h0408; // 0x1e84
	13'h0f43: q3 = 16'h8a04; // 0x1e86
	13'h0f44: q3 = 16'h0200; // 0x1e88
	13'h0f45: q3 = 16'h8a01; // 0x1e8a
	13'h0f46: q3 = 16'h0066; // 0x1e8c
	13'h0f47: q3 = 16'h8a08; // 0x1e8e
	13'h0f48: q3 = 16'h019a; // 0x1e90
	13'h0f49: q3 = 16'h8703; // 0x1e92
	13'h0f4a: q3 = 16'h0145; // 0x1e94
	13'h0f4b: q3 = 16'h03ce; // 0x1e96
	13'h0f4c: q3 = 16'h0400; // 0x1e98
	13'h0f4d: q3 = 16'h8a01; // 0x1e9a
	13'h0f4e: q3 = 16'h0400; // 0x1e9c
	13'h0f4f: q3 = 16'h8707; // 0x1e9e
	13'h0f50: q3 = 16'h016c; // 0x1ea0
	13'h0f51: q3 = 16'h0363; // 0x1ea2
	13'h0f52: q3 = 16'h088b; // 0x1ea4
	13'h0f53: q3 = 16'h0400; // 0x1ea6
	13'h0f54: q3 = 16'h8a05; // 0x1ea8
	13'h0f55: q3 = 16'h0400; // 0x1eaa
	13'h0f56: q3 = 16'h870f; // 0x1eac
	13'h0f57: q3 = 16'h0199; // 0x1eae
	13'h0f58: q3 = 16'h0333; // 0x1eb0
	13'h0f59: q3 = 16'h0666; // 0x1eb2
	13'h0f5a: q3 = 16'h0666; // 0x1eb4
	13'h0f5b: q3 = 16'h0400; // 0x1eb6
	13'h0f5c: q3 = 16'h8a01; // 0x1eb8
	13'h0f5d: q3 = 16'h0400; // 0x1eba
	13'h0f5e: q3 = 16'h0701; // 0x1ebc
	13'h0f5f: q3 = 16'h0222; // 0x1ebe
	13'h0f60: q3 = 16'h8a04; // 0x1ec0
	13'h0f61: q3 = 16'h0400; // 0x1ec2
	13'h0f62: q3 = 16'h8a01; // 0x1ec4
	13'h0f63: q3 = 16'h0266; // 0x1ec6
	13'h0f64: q3 = 16'h8a08; // 0x1ec8
	13'h0f65: q3 = 16'h019a; // 0x1eca
	13'h0f66: q3 = 16'h8703; // 0x1ecc
	13'h0f67: q3 = 16'h01e7; // 0x1ece
	13'h0f68: q3 = 16'h0445; // 0x1ed0
	13'h0f69: q3 = 16'h0400; // 0x1ed2
	13'h0f6a: q3 = 16'h8a01; // 0x1ed4
	13'h0f6b: q3 = 16'h0400; // 0x1ed6
	13'h0f6c: q3 = 16'h8701; // 0x1ed8
	13'h0f6d: q3 = 16'h01b1; // 0x1eda
	13'h0f6e: q3 = 16'h0400; // 0x1edc
	13'h0f6f: q3 = 16'h8a01; // 0x1ede
	13'h0f70: q3 = 16'h0400; // 0x1ee0
	13'h0f71: q3 = 16'h0302; // 0x1ee2
	13'h0f72: q3 = 16'h0000; // 0x1ee4
	13'h0f73: q3 = 16'hc314; // 0x1ee6
	13'h0f74: q3 = 16'h0502; // 0x1ee8
	13'h0f75: q3 = 16'h0000; // 0x1eea
	13'h0f76: q3 = 16'hc320; // 0x1eec
	13'h0f77: q3 = 16'h0a02; // 0x1eee
	13'h0f78: q3 = 16'h0100; // 0x1ef0
	13'h0f79: q3 = 16'hf667; // 0x1ef2
	13'h0f7a: q3 = 16'hf66b; // 0x1ef4
	13'h0f7b: q3 = 16'h000c; // 0x1ef6
	13'h0f7c: q3 = 16'h0700; // 0x1ef8
	13'h0f7d: q3 = 16'h0700; // 0x1efa
	13'h0f7e: q3 = 16'h0001; // 0x1efc
	13'h0f7f: q3 = 16'h0200; // 0x1efe
	13'h0f80: q3 = 16'h0200; // 0x1f00
	13'h0f81: q3 = 16'h0001; // 0x1f02
	13'h0f82: q3 = 16'hf980; // 0x1f04
	13'h0f83: q3 = 16'hf980; // 0x1f06
	13'h0f84: q3 = 16'h0002; // 0x1f08
	13'h0f85: q3 = 16'h04c0; // 0x1f0a
	13'h0f86: q3 = 16'h04c0; // 0x1f0c
	13'h0f87: q3 = 16'h0004; // 0x1f0e
	13'h0f88: q3 = 16'hfe29; // 0x1f10
	13'h0f89: q3 = 16'hfe2b; // 0x1f12
	13'h0f8a: q3 = 16'h0006; // 0x1f14
	13'h0f8b: q3 = 16'hfcaa; // 0x1f16
	13'h0f8c: q3 = 16'hfcab; // 0x1f18
	13'h0f8d: q3 = 16'h0003; // 0x1f1a
	13'h0f8e: q3 = 16'h0800; // 0x1f1c
	13'h0f8f: q3 = 16'h0800; // 0x1f1e
	13'h0f90: q3 = 16'h0002; // 0x1f20
	13'h0f91: q3 = 16'hfb40; // 0x1f22
	13'h0f92: q3 = 16'hfb40; // 0x1f24
	13'h0f93: q3 = 16'h0004; // 0x1f26
	13'h0f94: q3 = 16'hff80; // 0x1f28
	13'h0f95: q3 = 16'hff80; // 0x1f2a
	13'h0f96: q3 = 16'h0004; // 0x1f2c
	13'h0f97: q3 = 16'h0e00; // 0x1f2e
	13'h0f98: q3 = 16'h0e00; // 0x1f30
	13'h0f99: q3 = 16'h0002; // 0x1f32
	13'h0f9a: q3 = 16'hf400; // 0x1f34
	13'h0f9b: q3 = 16'hf400; // 0x1f36
	13'h0f9c: q3 = 16'h0002; // 0x1f38
	13'h0f9d: q3 = 16'hfd80; // 0x1f3a
	13'h0f9e: q3 = 16'hfd80; // 0x1f3c
	13'h0f9f: q3 = 16'h0002; // 0x1f3e
	13'h0fa0: q3 = 16'h0e00; // 0x1f40
	13'h0fa1: q3 = 16'h0e00; // 0x1f42
	13'h0fa2: q3 = 16'h0001; // 0x1f44
	13'h0fa3: q3 = 16'h0200; // 0x1f46
	13'h0fa4: q3 = 16'h0200; // 0x1f48
	13'h0fa5: q3 = 16'h0003; // 0x1f4a
	13'h0fa6: q3 = 16'hfbaa; // 0x1f4c
	13'h0fa7: q3 = 16'hfbab; // 0x1f4e
	13'h0fa8: q3 = 16'h0003; // 0x1f50
	13'h0fa9: q3 = 16'hfe40; // 0x1f52
	13'h0faa: q3 = 16'hfe40; // 0x1f54
	13'h0fab: q3 = 16'h0004; // 0x1f56
	13'h0fac: q3 = 16'h0000; // 0x1f58
	13'h0fad: q3 = 16'h0000; // 0x1f5a
	13'h0fae: q3 = 16'h0001; // 0x1f5c
	13'h0faf: q3 = 16'h0000; // 0x1f5e
	13'h0fb0: q3 = 16'h0000; // 0x1f60
	13'h0fb1: q3 = 16'h0001; // 0x1f62
	13'h0fb2: q3 = 16'h0200; // 0x1f64
	13'h0fb3: q3 = 16'h0200; // 0x1f66
	13'h0fb4: q3 = 16'h0002; // 0x1f68
	13'h0fb5: q3 = 16'hff00; // 0x1f6a
	13'h0fb6: q3 = 16'hff00; // 0x1f6c
	13'h0fb7: q3 = 16'h0004; // 0x1f6e
	13'h0fb8: q3 = 16'h0100; // 0x1f70
	13'h0fb9: q3 = 16'h0100; // 0x1f72
	13'h0fba: q3 = 16'h0001; // 0x1f74
	13'h0fbb: q3 = 16'h0600; // 0x1f76
	13'h0fbc: q3 = 16'h0600; // 0x1f78
	13'h0fbd: q3 = 16'h0001; // 0x1f7a
	13'h0fbe: q3 = 16'hfdaa; // 0x1f7c
	13'h0fbf: q3 = 16'hfdab; // 0x1f7e
	13'h0fc0: q3 = 16'h0003; // 0x1f80
	13'h0fc1: q3 = 16'h0800; // 0x1f82
	13'h0fc2: q3 = 16'h0800; // 0x1f84
	13'h0fc3: q3 = 16'h0002; // 0x1f86
	13'h0fc4: q3 = 16'h0000; // 0x1f88
	13'h0fc5: q3 = 16'h0000; // 0x1f8a
	13'h0fc6: q3 = 16'h0000; // 0x1f8c
	13'h0fc7: q3 = 16'h0097; // 0x1f8e
	13'h0fc8: q3 = 16'h0095; // 0x1f90
	13'h0fc9: q3 = 16'h0006; // 0x1f92
	13'h0fca: q3 = 16'h0008; // 0x1f94
	13'h0fcb: q3 = 16'h0005; // 0x1f96
	13'h0fcc: q3 = 16'h0019; // 0x1f98
	13'h0fcd: q3 = 16'h0000; // 0x1f9a
	13'h0fce: q3 = 16'h0000; // 0x1f9c
	13'h0fcf: q3 = 16'h0012; // 0x1f9e
	13'h0fd0: q3 = 16'hff20; // 0x1fa0
	13'h0fd1: q3 = 16'hff20; // 0x1fa2
	13'h0fd2: q3 = 16'h0004; // 0x1fa4
	13'h0fd3: q3 = 16'h0017; // 0x1fa6
	13'h0fd4: q3 = 16'h0015; // 0x1fa8
	13'h0fd5: q3 = 16'h0006; // 0x1faa
	13'h0fd6: q3 = 16'h0000; // 0x1fac
	13'h0fd7: q3 = 16'h0000; // 0x1fae
	13'h0fd8: q3 = 16'h0005; // 0x1fb0
	13'h0fd9: q3 = 16'h00c0; // 0x1fb2
	13'h0fda: q3 = 16'h00c0; // 0x1fb4
	13'h0fdb: q3 = 16'h0002; // 0x1fb6
	13'h0fdc: q3 = 16'h0000; // 0x1fb8
	13'h0fdd: q3 = 16'hf667; // 0x1fba
	13'h0fde: q3 = 16'h0000; // 0x1fbc
	13'h0fdf: q3 = 16'h00e0; // 0x1fbe
	13'h0fe0: q3 = 16'h0007; // 0x1fc0
	13'h0fe1: q3 = 16'h0000; // 0x1fc2
	13'h0fe2: q3 = 16'h0000; // 0x1fc4
	13'h0fe3: q3 = 16'h0000; // 0x1fc6
	13'h0fe4: q3 = 16'h8136; // 0x1fc8
	13'h0fe5: q3 = 16'h0000; // 0x1fca
	13'h0fe6: q3 = 16'hdef2; // 0x1fcc
	13'h0fe7: q3 = 16'h7f00; // 0x1fce
	13'h0fe8: q3 = 16'h0000; // 0x1fd0
	13'h0fe9: q3 = 16'h0000; // 0x1fd2
	13'h0fea: q3 = 16'h8136; // 0x1fd4
	13'h0feb: q3 = 16'h0000; // 0x1fd6
	13'h0fec: q3 = 16'hdf8e; // 0x1fd8
	13'h0fed: q3 = 16'h0000; // 0x1fda
	13'h0fee: q3 = 16'h0000; // 0x1fdc
	13'h0fef: q3 = 16'h0000; // 0x1fde
	13'h0ff0: q3 = 16'hdfbe; // 0x1fe0
	13'h0ff1: q3 = 16'h0000; // 0x1fe2
	13'h0ff2: q3 = 16'h0000; // 0x1fe4
	13'h0ff3: q3 = 16'h0514; // 0x1fe6
	13'h0ff4: q3 = 16'h0000; // 0x1fe8
	13'h0ff5: q3 = 16'h0000; // 0x1fea
	13'h0ff6: q3 = 16'hdfc6; // 0x1fec
	13'h0ff7: q3 = 16'hffff; // 0x1fee
	13'h0ff8: q3 = 16'h00b4; // 0x1ff0
	13'h0ff9: q3 = 16'h00aa; // 0x1ff2
	13'h0ffa: q3 = 16'h000f; // 0x1ff4
	13'h0ffb: q3 = 16'hfc00; // 0x1ff6
	13'h0ffc: q3 = 16'hfc00; // 0x1ff8
	13'h0ffd: q3 = 16'h0002; // 0x1ffa
	13'h0ffe: q3 = 16'h00c6; // 0x1ffc
	13'h0fff: q3 = 16'h00bb; // 0x1ffe
	13'h1000: q3 = 16'h000f; // 0x2000
	13'h1001: q3 = 16'hfb80; // 0x2002
	13'h1002: q3 = 16'hfb80; // 0x2004
	13'h1003: q3 = 16'h0002; // 0x2006
	13'h1004: q3 = 16'h00c0; // 0x2008
	13'h1005: q3 = 16'h00b4; // 0x200a
	13'h1006: q3 = 16'h0011; // 0x200c
	13'h1007: q3 = 16'hf700; // 0x200e
	13'h1008: q3 = 16'hf700; // 0x2010
	13'h1009: q3 = 16'h0001; // 0x2012
	13'h100a: q3 = 16'h0092; // 0x2014
	13'h100b: q3 = 16'h008e; // 0x2016
	13'h100c: q3 = 16'h0012; // 0x2018
	13'h100d: q3 = 16'hfa00; // 0x201a
	13'h100e: q3 = 16'hfa00; // 0x201c
	13'h100f: q3 = 16'h0001; // 0x201e
	13'h1010: q3 = 16'h0070; // 0x2020
	13'h1011: q3 = 16'h0069; // 0x2022
	13'h1012: q3 = 16'h0011; // 0x2024
	13'h1013: q3 = 16'h0000; // 0x2026
	13'h1014: q3 = 16'h0000; // 0x2028
	13'h1015: q3 = 16'h0000; // 0x202a
	13'h1016: q3 = 16'h03c0; // 0x202c
	13'h1017: q3 = 16'h03c0; // 0x202e
	13'h1018: q3 = 16'h0002; // 0x2030
	13'h1019: q3 = 16'hffce; // 0x2032
	13'h101a: q3 = 16'hffea; // 0x2034
	13'h101b: q3 = 16'h0056; // 0x2036
	13'h101c: q3 = 16'h0000; // 0x2038
	13'h101d: q3 = 16'h00b4; // 0x203a
	13'h101e: q3 = 16'h0000; // 0x203c
	13'h101f: q3 = 16'h0000; // 0x203e
	13'h1020: q3 = 16'h8136; // 0x2040
	13'h1021: q3 = 16'h0000; // 0x2042
	13'h1022: q3 = 16'hdff0; // 0x2044
	13'h1023: q3 = 16'h0600; // 0x2046
	13'h1024: q3 = 16'h0000; // 0x2048
	13'h1025: q3 = 16'h0000; // 0x204a
	13'h1026: q3 = 16'h8136; // 0x204c
	13'h1027: q3 = 16'h0000; // 0x204e
	13'h1028: q3 = 16'he02c; // 0x2050
	13'h1029: q3 = 16'h0000; // 0x2052
	13'h102a: q3 = 16'h0000; // 0x2054
	13'h102b: q3 = 16'h0000; // 0x2056
	13'h102c: q3 = 16'h0000; // 0x2058
	13'h102d: q3 = 16'h00e0; // 0x205a
	13'h102e: q3 = 16'h0000; // 0x205c
	13'h102f: q3 = 16'h05d2; // 0x205e
	13'h1030: q3 = 16'h0000; // 0x2060
	13'h1031: q3 = 16'h0000; // 0x2062
	13'h1032: q3 = 16'he03e; // 0x2064
	13'h1033: q3 = 16'hffff; // 0x2066
	13'h1034: q3 = 16'hffc6; // 0x2068
	13'h1035: q3 = 16'hffcd; // 0x206a
	13'h1036: q3 = 16'h0023; // 0x206c
	13'h1037: q3 = 16'h0600; // 0x206e
	13'h1038: q3 = 16'h0600; // 0x2070
	13'h1039: q3 = 16'h0001; // 0x2072
	13'h103a: q3 = 16'hffb4; // 0x2074
	13'h103b: q3 = 16'hffbb; // 0x2076
	13'h103c: q3 = 16'h0025; // 0x2078
	13'h103d: q3 = 16'h0900; // 0x207a
	13'h103e: q3 = 16'h0900; // 0x207c
	13'h103f: q3 = 16'h0001; // 0x207e
	13'h1040: q3 = 16'hff9a; // 0x2080
	13'h1041: q3 = 16'hffa6; // 0x2082
	13'h1042: q3 = 16'h0022; // 0x2084
	13'h1043: q3 = 16'h0240; // 0x2086
	13'h1044: q3 = 16'h0240; // 0x2088
	13'h1045: q3 = 16'h0004; // 0x208a
	13'h1046: q3 = 16'hff8c; // 0x208c
	13'h1047: q3 = 16'hffa6; // 0x208e
	13'h1048: q3 = 16'h001f; // 0x2090
	13'h1049: q3 = 16'h02ac; // 0x2092
	13'h104a: q3 = 16'h02aa; // 0x2094
	13'h104b: q3 = 16'h0003; // 0x2096
	13'h104c: q3 = 16'hff9c; // 0x2098
	13'h104d: q3 = 16'hffae; // 0x209a
	13'h104e: q3 = 16'h001f; // 0x209c
	13'h104f: q3 = 16'h0000; // 0x209e
	13'h1050: q3 = 16'h0000; // 0x20a0
	13'h1051: q3 = 16'h0000; // 0x20a2
	13'h1052: q3 = 16'h006b; // 0x20a4
	13'h1053: q3 = 16'h0009; // 0x20a6
	13'h1054: q3 = 16'h00ae; // 0x20a8
	13'h1055: q3 = 16'hfc40; // 0x20aa
	13'h1056: q3 = 16'hfc40; // 0x20ac
	13'h1057: q3 = 16'h0002; // 0x20ae
	13'h1058: q3 = 16'h0000; // 0x20b0
	13'h1059: q3 = 16'hffc6; // 0x20b2
	13'h105a: q3 = 16'h0000; // 0x20b4
	13'h105b: q3 = 16'h0000; // 0x20b6
	13'h105c: q3 = 16'h8136; // 0x20b8
	13'h105d: q3 = 16'h0000; // 0x20ba
	13'h105e: q3 = 16'he068; // 0x20bc
	13'h105f: q3 = 16'h1800; // 0x20be
	13'h1060: q3 = 16'h0000; // 0x20c0
	13'h1061: q3 = 16'h0000; // 0x20c2
	13'h1062: q3 = 16'h8136; // 0x20c4
	13'h1063: q3 = 16'h0000; // 0x20c6
	13'h1064: q3 = 16'he0a4; // 0x20c8
	13'h1065: q3 = 16'h0100; // 0x20ca
	13'h1066: q3 = 16'h0000; // 0x20cc
	13'h1067: q3 = 16'h0000; // 0x20ce
	13'h1068: q3 = 16'h0000; // 0x20d0
	13'h1069: q3 = 16'h00e0; // 0x20d2
	13'h106a: q3 = 16'h0000; // 0x20d4
	13'h106b: q3 = 16'h05dc; // 0x20d6
	13'h106c: q3 = 16'h0000; // 0x20d8
	13'h106d: q3 = 16'h0000; // 0x20da
	13'h106e: q3 = 16'he0b6; // 0x20dc
	13'h106f: q3 = 16'hffff; // 0x20de
	13'h1070: q3 = 16'h0000; // 0x20e0
	13'h1071: q3 = 16'h0006; // 0x20e2
	13'h1072: q3 = 16'h000d; // 0x20e4
	13'h1073: q3 = 16'h0011; // 0x20e6
	13'h1074: q3 = 16'h0015; // 0x20e8
	13'h1075: q3 = 16'h001b; // 0x20ea
	13'h1076: q3 = 16'h0024; // 0x20ec
	13'h1077: q3 = 16'h002b; // 0x20ee
	13'h1078: q3 = 16'h0031; // 0x20f0
	13'h1079: q3 = 16'h0039; // 0x20f2
	13'h107a: q3 = 16'h0045; // 0x20f4
	13'h107b: q3 = 16'h004d; // 0x20f6
	13'h107c: q3 = 16'h0054; // 0x20f8
	13'h107d: q3 = 16'h005d; // 0x20fa
	13'h107e: q3 = 16'h0066; // 0x20fc
	13'h107f: q3 = 16'h006b; // 0x20fe
	13'h1080: q3 = 16'h0071; // 0x2100
	13'h1081: q3 = 16'h0079; // 0x2102
	13'h1082: q3 = 16'h0083; // 0x2104
	13'h1083: q3 = 16'h008a; // 0x2106
	13'h1084: q3 = 16'h0091; // 0x2108
	13'h1085: q3 = 16'h009d; // 0x210a
	13'h1086: q3 = 16'h00a6; // 0x210c
	13'h1087: q3 = 16'h00ac; // 0x210e
	13'h1088: q3 = 16'h00b7; // 0x2110
	13'h1089: q3 = 16'h00c1; // 0x2112
	13'h108a: q3 = 16'h00ca; // 0x2114
	13'h108b: q3 = 16'h00ce; // 0x2116
	13'h108c: q3 = 16'h00d9; // 0x2118
	13'h108d: q3 = 16'h00e5; // 0x211a
	13'h108e: q3 = 16'h00f0; // 0x211c
	13'h108f: q3 = 16'h00f9; // 0x211e
	13'h1090: q3 = 16'h00fd; // 0x2120
	13'h1091: q3 = 16'h0108; // 0x2122
	13'h1092: q3 = 16'h0111; // 0x2124
	13'h1093: q3 = 16'h0116; // 0x2126
	13'h1094: q3 = 16'h0121; // 0x2128
	13'h1095: q3 = 16'h012f; // 0x212a
	13'h1096: q3 = 16'h0138; // 0x212c
	13'h1097: q3 = 16'h0140; // 0x212e
	13'h1098: q3 = 16'h014d; // 0x2130
	13'h1099: q3 = 16'h0152; // 0x2132
	13'h109a: q3 = 16'h0157; // 0x2134
	13'h109b: q3 = 16'h015c; // 0x2136
	13'h109c: q3 = 16'h0162; // 0x2138
	13'h109d: q3 = 16'h0179; // 0x213a
	13'h109e: q3 = 16'h018b; // 0x213c
	13'h109f: q3 = 16'h01a3; // 0x213e
	13'h10a0: q3 = 16'h01bc; // 0x2140
	13'h10a1: q3 = 16'h01bd; // 0x2142
	13'h10a2: q3 = 16'h01cc; // 0x2144
	13'h10a3: q3 = 16'h01e4; // 0x2146
	13'h10a4: q3 = 16'h01ec; // 0x2148
	13'h10a5: q3 = 16'h01fe; // 0x214a
	13'h10a6: q3 = 16'h0213; // 0x214c
	13'h10a7: q3 = 16'h022a; // 0x214e
	13'h10a8: q3 = 16'h0241; // 0x2150
	13'h10a9: q3 = 16'h0246; // 0x2152
	13'h10aa: q3 = 16'h024b; // 0x2154
	13'h10ab: q3 = 16'h0253; // 0x2156
	13'h10ac: q3 = 16'h0259; // 0x2158
	13'h10ad: q3 = 16'h0268; // 0x215a
	13'h10ae: q3 = 16'h0277; // 0x215c
	13'h10af: q3 = 16'h0289; // 0x215e
	13'h10b0: q3 = 16'h029f; // 0x2160
	13'h10b1: q3 = 16'h02a2; // 0x2162
	13'h10b2: q3 = 16'h02a6; // 0x2164
	13'h10b3: q3 = 16'h02ac; // 0x2166
	13'h10b4: q3 = 16'h02af; // 0x2168
	13'h10b5: q3 = 16'h02b7; // 0x216a
	13'h10b6: q3 = 16'h02ba; // 0x216c
	13'h10b7: q3 = 16'h02c2; // 0x216e
	13'h10b8: q3 = 16'h02ca; // 0x2170
	13'h10b9: q3 = 16'h02ce; // 0x2172
	13'h10ba: q3 = 16'h02d2; // 0x2174
	13'h10bb: q3 = 16'h02d5; // 0x2176
	13'h10bc: q3 = 16'h02d8; // 0x2178
	13'h10bd: q3 = 16'h02df; // 0x217a
	13'h10be: q3 = 16'h02e8; // 0x217c
	13'h10bf: q3 = 16'h02f5; // 0x217e
	13'h10c0: q3 = 16'h0300; // 0x2180
	13'h10c1: q3 = 16'h0308; // 0x2182
	13'h10c2: q3 = 16'h030b; // 0x2184
	13'h10c3: q3 = 16'h0313; // 0x2186
	13'h10c4: q3 = 16'h0316; // 0x2188
	13'h10c5: q3 = 16'h031a; // 0x218a
	13'h10c6: q3 = 16'h031e; // 0x218c
	13'h10c7: q3 = 16'h0321; // 0x218e
	13'h10c8: q3 = 16'h0328; // 0x2190
	13'h10c9: q3 = 16'h033d; // 0x2192
	13'h10ca: q3 = 16'h0352; // 0x2194
	13'h10cb: q3 = 16'h0367; // 0x2196
	13'h10cc: q3 = 16'h037d; // 0x2198
	13'h10cd: q3 = 16'h0389; // 0x219a
	13'h10ce: q3 = 16'h0398; // 0x219c
	13'h10cf: q3 = 16'h03a4; // 0x219e
	13'h10d0: q3 = 16'h03af; // 0x21a0
	13'h10d1: q3 = 16'h03b8; // 0x21a2
	13'h10d2: q3 = 16'h03c8; // 0x21a4
	13'h10d3: q3 = 16'h03d7; // 0x21a6
	13'h10d4: q3 = 16'h03e0; // 0x21a8
	13'h10d5: q3 = 16'h03f0; // 0x21aa
	13'h10d6: q3 = 16'h03fe; // 0x21ac
	13'h10d7: q3 = 16'h0416; // 0x21ae
	13'h10d8: q3 = 16'h0427; // 0x21b0
	13'h10d9: q3 = 16'h0428; // 0x21b2
	13'h10da: q3 = 16'h0429; // 0x21b4
	13'h10db: q3 = 16'h0436; // 0x21b6
	13'h10dc: q3 = 16'h0442; // 0x21b8
	13'h10dd: q3 = 16'h0458; // 0x21ba
	13'h10de: q3 = 16'h046d; // 0x21bc
	13'h10df: q3 = 16'h047e; // 0x21be
	13'h10e0: q3 = 16'h048d; // 0x21c0
	13'h10e1: q3 = 16'h049c; // 0x21c2
	13'h10e2: q3 = 16'h04ab; // 0x21c4
	13'h10e3: q3 = 16'h04c3; // 0x21c6
	13'h10e4: q3 = 16'h04d2; // 0x21c8
	13'h10e5: q3 = 16'h04e4; // 0x21ca
	13'h10e6: q3 = 16'h04f8; // 0x21cc
	13'h10e7: q3 = 16'h0511; // 0x21ce
	13'h10e8: q3 = 16'h0527; // 0x21d0
	13'h10e9: q3 = 16'h0528; // 0x21d2
	13'h10ea: q3 = 16'h0529; // 0x21d4
	13'h10eb: q3 = 16'h053b; // 0x21d6
	13'h10ec: q3 = 16'h053c; // 0x21d8
	13'h10ed: q3 = 16'h054b; // 0x21da
	13'h10ee: q3 = 16'h055d; // 0x21dc
	13'h10ef: q3 = 16'h056f; // 0x21de
	13'h10f0: q3 = 16'h0587; // 0x21e0
	13'h10f1: q3 = 16'h0593; // 0x21e2
	13'h10f2: q3 = 16'h059f; // 0x21e4
	13'h10f3: q3 = 16'h05b3; // 0x21e6
	13'h10f4: q3 = 16'h05cb; // 0x21e8
	13'h10f5: q3 = 16'h05dd; // 0x21ea
	13'h10f6: q3 = 16'h05e5; // 0x21ec
	13'h10f7: q3 = 16'h05fe; // 0x21ee
	13'h10f8: q3 = 16'h0611; // 0x21f0
	13'h10f9: q3 = 16'h0618; // 0x21f2
	13'h10fa: q3 = 16'h0624; // 0x21f4
	13'h10fb: q3 = 16'h0637; // 0x21f6
	13'h10fc: q3 = 16'h063e; // 0x21f8
	13'h10fd: q3 = 16'h0653; // 0x21fa
	13'h10fe: q3 = 16'h0663; // 0x21fc
	13'h10ff: q3 = 16'h0672; // 0x21fe
	13'h1100: q3 = 16'h067e; // 0x2200
	13'h1101: q3 = 16'h067f; // 0x2202
	13'h1102: q3 = 16'h068b; // 0x2204
	13'h1103: q3 = 16'h069c; // 0x2206
	13'h1104: q3 = 16'h06a9; // 0x2208
	13'h1105: q3 = 16'h06b9; // 0x220a
	13'h1106: q3 = 16'h06c9; // 0x220c
	13'h1107: q3 = 16'h06de; // 0x220e
	13'h1108: q3 = 16'h06f4; // 0x2210
	13'h1109: q3 = 16'h06fd; // 0x2212
	13'h110a: q3 = 16'h0706; // 0x2214
	13'h110b: q3 = 16'h071f; // 0x2216
	13'h110c: q3 = 16'h0734; // 0x2218
	13'h110d: q3 = 16'h0735; // 0x221a
	13'h110e: q3 = 16'h0736; // 0x221c
	13'h110f: q3 = 16'h073f; // 0x221e
	13'h1110: q3 = 16'h0740; // 0x2220
	13'h1111: q3 = 16'h0753; // 0x2222
	13'h1112: q3 = 16'h0766; // 0x2224
	13'h1113: q3 = 16'h0777; // 0x2226
	13'h1114: q3 = 16'h078c; // 0x2228
	13'h1115: q3 = 16'h0793; // 0x222a
	13'h1116: q3 = 16'h0799; // 0x222c
	13'h1117: q3 = 16'h07a0; // 0x222e
	13'h1118: q3 = 16'h07a7; // 0x2230
	13'h1119: q3 = 16'h07ae; // 0x2232
	13'h111a: q3 = 16'h07b4; // 0x2234
	13'h111b: q3 = 16'h07bb; // 0x2236
	13'h111c: q3 = 16'h07c2; // 0x2238
	13'h111d: q3 = 16'h07d2; // 0x223a
	13'h111e: q3 = 16'h07e5; // 0x223c
	13'h111f: q3 = 16'h07fb; // 0x223e
	13'h1120: q3 = 16'h0811; // 0x2240
	13'h1121: q3 = 16'h0826; // 0x2242
	13'h1122: q3 = 16'h083a; // 0x2244
	13'h1123: q3 = 16'h0845; // 0x2246
	13'h1124: q3 = 16'h084f; // 0x2248
	13'h1125: q3 = 16'h0858; // 0x224a
	13'h1126: q3 = 16'h0865; // 0x224c
	13'h1127: q3 = 16'h0871; // 0x224e
	13'h1128: q3 = 16'h087f; // 0x2250
	13'h1129: q3 = 16'h088d; // 0x2252
	13'h112a: q3 = 16'h089c; // 0x2254
	13'h112b: q3 = 16'h08b1; // 0x2256
	13'h112c: q3 = 16'h08c4; // 0x2258
	13'h112d: q3 = 16'h08c8; // 0x225a
	13'h112e: q3 = 16'h08cd; // 0x225c
	13'h112f: q3 = 16'h08d3; // 0x225e
	13'h1130: q3 = 16'h08d9; // 0x2260
	13'h1131: q3 = 16'h08df; // 0x2262
	13'h1132: q3 = 16'h08e8; // 0x2264
	13'h1133: q3 = 16'h08ee; // 0x2266
	13'h1134: q3 = 16'h08f3; // 0x2268
	13'h1135: q3 = 16'h0908; // 0x226a
	13'h1136: q3 = 16'h0920; // 0x226c
	13'h1137: q3 = 16'h092f; // 0x226e
	13'h1138: q3 = 16'h093e; // 0x2270
	13'h1139: q3 = 16'h093f; // 0x2272
	13'h113a: q3 = 16'h0940; // 0x2274
	13'h113b: q3 = 16'h094c; // 0x2276
	13'h113c: q3 = 16'h095b; // 0x2278
	13'h113d: q3 = 16'h096a; // 0x227a
	13'h113e: q3 = 16'h097b; // 0x227c
	13'h113f: q3 = 16'h0993; // 0x227e
	13'h1140: q3 = 16'h09a5; // 0x2280
	13'h1141: q3 = 16'h09b7; // 0x2282
	13'h1142: q3 = 16'h09c3; // 0x2284
	13'h1143: q3 = 16'h09d4; // 0x2286
	13'h1144: q3 = 16'h09e8; // 0x2288
	13'h1145: q3 = 16'h09f4; // 0x228a
	13'h1146: q3 = 16'h09fe; // 0x228c
	13'h1147: q3 = 16'h0a10; // 0x228e
	13'h1148: q3 = 16'h0a22; // 0x2290
	13'h1149: q3 = 16'h0a2e; // 0x2292
	13'h114a: q3 = 16'h0a3a; // 0x2294
	13'h114b: q3 = 16'h0a4c; // 0x2296
	13'h114c: q3 = 16'h0a5b; // 0x2298
	13'h114d: q3 = 16'h0a61; // 0x229a
	13'h114e: q3 = 16'h0a68; // 0x229c
	13'h114f: q3 = 16'h0a6f; // 0x229e
	13'h1150: q3 = 16'h0a75; // 0x22a0
	13'h1151: q3 = 16'h0a7b; // 0x22a2
	13'h1152: q3 = 16'h0a81; // 0x22a4
	13'h1153: q3 = 16'h0a88; // 0x22a6
	13'h1154: q3 = 16'h0a8e; // 0x22a8
	13'h1155: q3 = 16'h0a92; // 0x22aa
	13'h1156: q3 = 16'h0a99; // 0x22ac
	13'h1157: q3 = 16'h0aa0; // 0x22ae
	13'h1158: q3 = 16'h0aa6; // 0x22b0
	13'h1159: q3 = 16'h0aaa; // 0x22b2
	13'h115a: q3 = 16'h0ab0; // 0x22b4
	13'h115b: q3 = 16'h0ab8; // 0x22b6
	13'h115c: q3 = 16'h0abc; // 0x22b8
	13'h115d: q3 = 16'h0ac3; // 0x22ba
	13'h115e: q3 = 16'h0ac9; // 0x22bc
	13'h115f: q3 = 16'h0acf; // 0x22be
	13'h1160: q3 = 16'h0ad5; // 0x22c0
	13'h1161: q3 = 16'h0ade; // 0x22c2
	13'h1162: q3 = 16'h0ae8; // 0x22c4
	13'h1163: q3 = 16'h0aee; // 0x22c6
	13'h1164: q3 = 16'h0af5; // 0x22c8
	13'h1165: q3 = 16'h0b0e; // 0x22ca
	13'h1166: q3 = 16'h0b10; // 0x22cc
	13'h1167: q3 = 16'h0b1c; // 0x22ce
	13'h1168: q3 = 16'h0b25; // 0x22d0
	13'h1169: q3 = 16'h0b2e; // 0x22d2
	13'h116a: q3 = 16'h0b34; // 0x22d4
	13'h116b: q3 = 16'h0b3d; // 0x22d6
	13'h116c: q3 = 16'h0b43; // 0x22d8
	13'h116d: q3 = 16'h0b48; // 0x22da
	13'h116e: q3 = 16'h0b4e; // 0x22dc
	13'h116f: q3 = 16'h0b53; // 0x22de
	13'h1170: q3 = 16'h0b58; // 0x22e0
	13'h1171: q3 = 16'h0b5e; // 0x22e2
	13'h1172: q3 = 16'h0b6b; // 0x22e4
	13'h1173: q3 = 16'h0b77; // 0x22e6
	13'h1174: q3 = 16'h0b85; // 0x22e8
	13'h1175: q3 = 16'h0b94; // 0x22ea
	13'h1176: q3 = 16'h0b9a; // 0x22ec
	13'h1177: q3 = 16'h0bab; // 0x22ee
	13'h1178: q3 = 16'h0bb5; // 0x22f0
	13'h1179: q3 = 16'h0bc2; // 0x22f2
	13'h117a: q3 = 16'h0bca; // 0x22f4
	13'h117b: q3 = 16'h0bd2; // 0x22f6
	13'h117c: q3 = 16'h0bdd; // 0x22f8
	13'h117d: q3 = 16'h0be7; // 0x22fa
	13'h117e: q3 = 16'h0be9; // 0x22fc
	13'h117f: q3 = 16'h0bf2; // 0x22fe
	13'h1180: q3 = 16'h0c07; // 0x2300
	13'h1181: q3 = 16'h0c0c; // 0x2302
	13'h1182: q3 = 16'h0c15; // 0x2304
	13'h1183: q3 = 16'h0c1b; // 0x2306
	13'h1184: q3 = 16'h0c23; // 0x2308
	13'h1185: q3 = 16'h0c35; // 0x230a
	13'h1186: q3 = 16'h0c45; // 0x230c
	13'h1187: q3 = 16'h0c5e; // 0x230e
	13'h1188: q3 = 16'h0c6e; // 0x2310
	13'h1189: q3 = 16'h0c77; // 0x2312
	13'h118a: q3 = 16'h0c82; // 0x2314
	13'h118b: q3 = 16'h0c91; // 0x2316
	13'h118c: q3 = 16'h0c9a; // 0x2318
	13'h118d: q3 = 16'h0c9f; // 0x231a
	13'h118e: q3 = 16'h0cb3; // 0x231c
	13'h118f: q3 = 16'h0cc3; // 0x231e
	13'h1190: q3 = 16'h0cdb; // 0x2320
	13'h1191: q3 = 16'h0ce8; // 0x2322
	13'h1192: q3 = 16'h0cfc; // 0x2324
	13'h1193: q3 = 16'h0d0a; // 0x2326
	13'h1194: q3 = 16'h0d19; // 0x2328
	13'h1195: q3 = 16'h0d22; // 0x232a
	13'h1196: q3 = 16'h0d2b; // 0x232c
	13'h1197: q3 = 16'h0d3a; // 0x232e
	13'h1198: q3 = 16'h0d43; // 0x2330
	13'h1199: q3 = 16'h0d5b; // 0x2332
	13'h119a: q3 = 16'h0d61; // 0x2334
	13'h119b: q3 = 16'h0d67; // 0x2336
	13'h119c: q3 = 16'h0d6d; // 0x2338
	13'h119d: q3 = 16'h0d76; // 0x233a
	13'h119e: q3 = 16'h0d79; // 0x233c
	13'h119f: q3 = 16'h0d7c; // 0x233e
	13'h11a0: q3 = 16'h0d84; // 0x2340
	13'h11a1: q3 = 16'h0d8d; // 0x2342
	13'h11a2: q3 = 16'h0d94; // 0x2344
	13'h11a3: q3 = 16'h0dac; // 0x2346
	13'h11a4: q3 = 16'h0db2; // 0x2348
	13'h11a5: q3 = 16'h0dbb; // 0x234a
	13'h11a6: q3 = 16'h0dbe; // 0x234c
	13'h11a7: q3 = 16'h0dc1; // 0x234e
	13'h11a8: q3 = 16'h0dc7; // 0x2350
	13'h11a9: q3 = 16'h0ddc; // 0x2352
	13'h11aa: q3 = 16'h0df3; // 0x2354
	13'h11ab: q3 = 16'h0e02; // 0x2356
	13'h11ac: q3 = 16'h0e09; // 0x2358
	13'h11ad: q3 = 16'h0e16; // 0x235a
	13'h11ae: q3 = 16'h0e20; // 0x235c
	13'h11af: q3 = 16'h0e2c; // 0x235e
	13'h11b0: q3 = 16'h0e35; // 0x2360
	13'h11b1: q3 = 16'h0e43; // 0x2362
	13'h11b2: q3 = 16'h0e52; // 0x2364
	13'h11b3: q3 = 16'h0e61; // 0x2366
	13'h11b4: q3 = 16'h0e6f; // 0x2368
	13'h11b5: q3 = 16'h0e7b; // 0x236a
	13'h11b6: q3 = 16'h0e82; // 0x236c
	13'h11b7: q3 = 16'h0e8d; // 0x236e
	13'h11b8: q3 = 16'h0e98; // 0x2370
	13'h11b9: q3 = 16'h0e9e; // 0x2372
	13'h11ba: q3 = 16'h0ea4; // 0x2374
	13'h11bb: q3 = 16'h0ead; // 0x2376
	13'h11bc: q3 = 16'h0eb6; // 0x2378
	13'h11bd: q3 = 16'h0eb8; // 0x237a
	13'h11be: q3 = 16'h0eba; // 0x237c
	13'h11bf: q3 = 16'h0ebc; // 0x237e
	13'h11c0: q3 = 16'h0ebe; // 0x2380
	13'h11c1: q3 = 16'h0ec0; // 0x2382
	13'h11c2: q3 = 16'h0ec3; // 0x2384
	13'h11c3: q3 = 16'h0ec6; // 0x2386
	13'h11c4: q3 = 16'h0ecc; // 0x2388
	13'h11c5: q3 = 16'h0ed3; // 0x238a
	13'h11c6: q3 = 16'h0ed7; // 0x238c
	13'h11c7: q3 = 16'h0eda; // 0x238e
	13'h11c8: q3 = 16'h0ee0; // 0x2390
	13'h11c9: q3 = 16'h0ee6; // 0x2392
	13'h11ca: q3 = 16'h0eec; // 0x2394
	13'h11cb: q3 = 16'h0ef2; // 0x2396
	13'h11cc: q3 = 16'h0ef5; // 0x2398
	13'h11cd: q3 = 16'h0ef8; // 0x239a
	13'h11ce: q3 = 16'h0efa; // 0x239c
	13'h11cf: q3 = 16'h0f03; // 0x239e
	13'h11d0: q3 = 16'h0f0a; // 0x23a0
	13'h11d1: q3 = 16'h0f0c; // 0x23a2
	13'h11d2: q3 = 16'h0f15; // 0x23a4
	13'h11d3: q3 = 16'h0f1b; // 0x23a6
	13'h11d4: q3 = 16'h0f24; // 0x23a8
	13'h11d5: q3 = 16'h0f30; // 0x23aa
	13'h11d6: q3 = 16'h0f39; // 0x23ac
	13'h11d7: q3 = 16'h0f3f; // 0x23ae
	13'h11d8: q3 = 16'h0f4b; // 0x23b0
	13'h11d9: q3 = 16'h0f56; // 0x23b2
	13'h11da: q3 = 16'h0000; // 0x23b4
	13'h11db: q3 = 16'hff00; // 0x23b6
	13'h11dc: q3 = 16'h8ef9; // 0x23b8
	13'h11dd: q3 = 16'ha696; // 0x23ba
	13'h11de: q3 = 16'h5f80; // 0x23bc
	13'h11df: q3 = 16'hae19; // 0x23be
	13'h11e0: q3 = 16'ha696; // 0x23c0
	13'h11e1: q3 = 16'h5a73; // 0x23c2
	13'h11e2: q3 = 16'hf88e; // 0x23c4
	13'h11e3: q3 = 16'h19a5; // 0x23c6
	13'h11e4: q3 = 16'hf88e; // 0x23c8
	13'h11e5: q3 = 16'h19a5; // 0x23ca
	13'h11e6: q3 = 16'hf8da; // 0x23cc
	13'h11e7: q3 = 16'h1ba9; // 0x23ce
	13'h11e8: q3 = 16'hb2c8; // 0x23d0
	13'h11e9: q3 = 16'h7eda; // 0x23d2
	13'h11ea: q3 = 16'h1ba9; // 0x23d4
	13'h11eb: q3 = 16'hb2c9; // 0x23d6
	13'h11ec: q3 = 16'h65a7; // 0x23d8
	13'h11ed: q3 = 16'h3f80; // 0x23da
	13'h11ee: q3 = 16'hda1a; // 0x23dc
	13'h11ef: q3 = 16'h6ea6; // 0x23de
	13'h11f0: q3 = 16'hcb21; // 0x23e0
	13'h11f1: q3 = 16'hf8da; // 0x23e2
	13'h11f2: q3 = 16'h1ba9; // 0x23e4
	13'h11f3: q3 = 16'hb2c9; // 0x23e6
	13'h11f4: q3 = 16'h7e8e; // 0x23e8
	13'h11f5: q3 = 16'h8be3; // 0x23ea
	13'h11f6: q3 = 16'hbec8; // 0x23ec
	13'h11f7: q3 = 16'h7497; // 0x23ee
	13'h11f8: q3 = 16'he0ce; // 0x23f0
	13'h11f9: q3 = 16'h3a2f; // 0x23f2
	13'h11fa: q3 = 16'haefb; // 0x23f4
	13'h11fb: q3 = 16'h2192; // 0x23f6
	13'h11fc: q3 = 16'h5ba5; // 0x23f8
	13'h11fd: q3 = 16'ha73f; // 0x23fa
	13'h11fe: q3 = 16'h808e; // 0x23fc
	13'h11ff: q3 = 16'h8be3; // 0x23fe
	13'h1200: q3 = 16'hbec8; // 0x2400
	13'h1201: q3 = 16'h7497; // 0x2402
	13'h1202: q3 = 16'he08e; // 0x2404
	13'h1203: q3 = 16'h8be3; // 0x2406
	13'h1204: q3 = 16'hbec8; // 0x2408
	13'h1205: q3 = 16'h74f8; // 0x240a
	13'h1206: q3 = 16'hcf4c; // 0x240c
	13'h1207: q3 = 16'ha1de; // 0x240e
	13'h1208: q3 = 16'h2972; // 0x2410
	13'h1209: q3 = 16'hcb9f; // 0x2412
	13'h120a: q3 = 16'h8097; // 0x2414
	13'h120b: q3 = 16'h2922; // 0x2416
	13'h120c: q3 = 16'h965c; // 0x2418
	13'h120d: q3 = 16'ha5a7; // 0x241a
	13'h120e: q3 = 16'h3f80; // 0x241c
	13'h120f: q3 = 16'h9b29; // 0x241e
	13'h1210: q3 = 16'h7387; // 0x2420
	13'h1211: q3 = 16'he09b; // 0x2422
	13'h1212: q3 = 16'h2869; // 0x2424
	13'h1213: q3 = 16'hce5f; // 0x2426
	13'h1214: q3 = 16'h80c2; // 0x2428
	13'h1215: q3 = 16'h9cf4; // 0x242a
	13'h1216: q3 = 16'h863a; // 0x242c
	13'h1217: q3 = 16'h29bf; // 0x242e
	13'h1218: q3 = 16'he0c2; // 0x2430
	13'h1219: q3 = 16'h9cf4; // 0x2432
	13'h121a: q3 = 16'h87aa; // 0x2434
	13'h121b: q3 = 16'h65ba; // 0x2436
	13'h121c: q3 = 16'h5a73; // 0x2438
	13'h121d: q3 = 16'hf8c2; // 0x243a
	13'h121e: q3 = 16'h9cf4; // 0x243c
	13'h121f: q3 = 16'h863a; // 0x243e
	13'h1220: q3 = 16'h2ff8; // 0x2440
	13'h1221: q3 = 16'hc29c; // 0x2442
	13'h1222: q3 = 16'hf486; // 0x2444
	13'h1223: q3 = 16'h3a25; // 0x2446
	13'h1224: q3 = 16'hf8bf; // 0x2448
	13'h1225: q3 = 16'h286e; // 0x244a
	13'h1226: q3 = 16'h9e50; // 0x244c
	13'h1227: q3 = 16'h33a2; // 0x244e
	13'h1228: q3 = 16'h5ca2; // 0x2450
	13'h1229: q3 = 16'h974f; // 0x2452
	13'h122a: q3 = 16'h80bf; // 0x2454
	13'h122b: q3 = 16'h286e; // 0x2456
	13'h122c: q3 = 16'h9e5b; // 0x2458
	13'h122d: q3 = 16'ha5a7; // 0x245a
	13'h122e: q3 = 16'h3f80; // 0x245c
	13'h122f: q3 = 16'hba1c; // 0x245e
	13'h1230: q3 = 16'ha1ba; // 0x2460
	13'h1231: q3 = 16'ha87e; // 0x2462
	13'h1232: q3 = 16'hcefc; // 0x2464
	13'h1233: q3 = 16'ha297; // 0x2466
	13'h1234: q3 = 16'h402f; // 0x2468
	13'h1235: q3 = 16'hca1b; // 0x246a
	13'h1236: q3 = 16'ha797; // 0x246c
	13'h1237: q3 = 16'he0b2; // 0x246e
	13'h1238: q3 = 16'h9b65; // 0x2470
	13'h1239: q3 = 16'h033a; // 0x2472
	13'h123a: q3 = 16'h25ca; // 0x2474
	13'h123b: q3 = 16'h2974; // 0x2476
	13'h123c: q3 = 16'hf8b2; // 0x2478
	13'h123d: q3 = 16'h9b6f; // 0x247a
	13'h123e: q3 = 16'hba5b; // 0x247c
	13'h123f: q3 = 16'ha5a7; // 0x247e
	13'h1240: q3 = 16'h3f80; // 0x2480
	13'h1241: q3 = 16'hb29b; // 0x2482
	13'h1242: q3 = 16'h61f8; // 0x2484
	13'h1243: q3 = 16'hcefc; // 0x2486
	13'h1244: q3 = 16'ha297; // 0x2488
	13'h1245: q3 = 16'h402d; // 0x248a
	13'h1246: q3 = 16'h96ed; // 0x248c
	13'h1247: q3 = 16'h2897; // 0x248e
	13'h1248: q3 = 16'he08a; // 0x2490
	13'h1249: q3 = 16'hc863; // 0x2492
	13'h124a: q3 = 16'hac0c; // 0x2494
	13'h124b: q3 = 16'ha1cf; // 0x2496
	13'h124c: q3 = 16'h08a5; // 0x2498
	13'h124d: q3 = 16'hcb2e; // 0x249a
	13'h124e: q3 = 16'h7e8b; // 0x249c
	13'h124f: q3 = 16'h2bed; // 0x249e
	13'h1250: q3 = 16'h8a59; // 0x24a0
	13'h1251: q3 = 16'h7296; // 0x24a2
	13'h1252: q3 = 16'he969; // 0x24a4
	13'h1253: q3 = 16'hcfe0; // 0x24a6
	13'h1254: q3 = 16'hb6fc; // 0x24a8
	13'h1255: q3 = 16'ha102; // 0x24aa
	13'h1256: q3 = 16'he967; // 0x24ac
	13'h1257: q3 = 16'hca1f; // 0x24ae
	13'h1258: q3 = 16'h80b7; // 0x24b0
	13'h1259: q3 = 16'h5ca5; // 0x24b2
	13'h125a: q3 = 16'hf8b2; // 0x24b4
	13'h125b: q3 = 16'h5b6f; // 0x24b6
	13'h125c: q3 = 16'hb80c; // 0x24b8
	13'h125d: q3 = 16'he897; // 0x24ba
	13'h125e: q3 = 16'h28a5; // 0x24bc
	13'h125f: q3 = 16'hd3e0; // 0x24be
	13'h1260: q3 = 16'hea9d; // 0x24c0
	13'h1261: q3 = 16'h32be; // 0x24c2
	13'h1262: q3 = 16'he96e; // 0x24c4
	13'h1263: q3 = 16'h969c; // 0x24c6
	13'h1264: q3 = 16'hfeb2; // 0x24c8
	13'h1265: q3 = 16'h9b6f; // 0x24ca
	13'h1266: q3 = 16'hbbe0; // 0x24cc
	13'h1267: q3 = 16'hcefc; // 0x24ce
	13'h1268: q3 = 16'ha297; // 0x24d0
	13'h1269: q3 = 16'h4023; // 0x24d2
	13'h126a: q3 = 16'ha74c; // 0x24d4
	13'h126b: q3 = 16'hafbb; // 0x24d6
	13'h126c: q3 = 16'he0ca; // 0x24d8
	13'h126d: q3 = 16'h1cf0; // 0x24da
	13'h126e: q3 = 16'h8a5c; // 0x24dc
	13'h126f: q3 = 16'hb2e4; // 0x24de
	13'h1270: q3 = 16'h0ce8; // 0x24e0
	13'h1271: q3 = 16'h9728; // 0x24e2
	13'h1272: q3 = 16'ha5d3; // 0x24e4
	13'h1273: q3 = 16'he0a2; // 0x24e6
	13'h1274: q3 = 16'h9b62; // 0x24e8
	13'h1275: q3 = 16'h965c; // 0x24ea
	13'h1276: q3 = 16'ha5a7; // 0x24ec
	13'h1277: q3 = 16'h3f80; // 0x24ee
	13'h1278: q3 = 16'h9b28; // 0x24f0
	13'h1279: q3 = 16'h6d8b; // 0x24f2
	13'h127a: q3 = 16'h5973; // 0x24f4
	13'h127b: q3 = 16'h87e0; // 0x24f6
	13'h127c: q3 = 16'hcefc; // 0x24f8
	13'h127d: q3 = 16'ha297; // 0x24fa
	13'h127e: q3 = 16'h4026; // 0x24fc
	13'h127f: q3 = 16'hca1b; // 0x24fe
	13'h1280: q3 = 16'h62be; // 0x2500
	13'h1281: q3 = 16'h9ce5; // 0x2502
	13'h1282: q3 = 16'hf8b2; // 0x2504
	13'h1283: q3 = 16'h5da5; // 0x2506
	13'h1284: q3 = 16'hb3e0; // 0x2508
	13'h1285: q3 = 16'hcf4d; // 0x250a
	13'h1286: q3 = 16'h6697; // 0x250c
	13'h1287: q3 = 16'he0ba; // 0x250e
	13'h1288: q3 = 16'h9da5; // 0x2510
	13'h1289: q3 = 16'hb3e0; // 0x2512
	13'h128a: q3 = 16'hba9d; // 0x2514
	13'h128b: q3 = 16'ha587; // 0x2516
	13'h128c: q3 = 16'h5f80; // 0x2518
	13'h128d: q3 = 16'hb6fd; // 0x251a
	13'h128e: q3 = 16'ha502; // 0x251c
	13'h128f: q3 = 16'habf9; // 0x251e
	13'h1290: q3 = 16'hcf4a; // 0x2520
	13'h1291: q3 = 16'h63ac; // 0x2522
	13'h1292: q3 = 16'h0d2f; // 0x2524
	13'h1293: q3 = 16'h0339; // 0x2526
	13'h1294: q3 = 16'h6c96; // 0x2528
	13'h1295: q3 = 16'h3d00; // 0x252a
	13'h1296: q3 = 16'hb25d; // 0x252c
	13'h1297: q3 = 16'ha5b3; // 0x252e
	13'h1298: q3 = 16'he0cf; // 0x2530
	13'h1299: q3 = 16'h4975; // 0x2532
	13'h129a: q3 = 16'h972a; // 0x2534
	13'h129b: q3 = 16'heed6; // 0x2536
	13'h129c: q3 = 16'h5c30; // 0x2538
	13'h129d: q3 = 16'h96c0; // 0x253a
	13'h129e: q3 = 16'h2297; // 0x253c
	13'h129f: q3 = 16'h7967; // 0x253e
	13'h12a0: q3 = 16'h96e3; // 0x2540
	13'h12a1: q3 = 16'h3eb6; // 0x2542
	13'h12a2: q3 = 16'hfda5; // 0x2544
	13'h12a3: q3 = 16'hc80b; // 0x2546
	13'h12a4: q3 = 16'h2103; // 0x2548
	13'h12a5: q3 = 16'h086c; // 0x254a
	13'h12a6: q3 = 16'h86e8; // 0x254c
	13'h12a7: q3 = 16'he102; // 0x254e
	13'h12a8: q3 = 16'h4940; // 0x2550
	13'h12a9: q3 = 16'hb61b; // 0x2552
	13'h12aa: q3 = 16'ha4bc; // 0x2554
	13'h12ab: q3 = 16'h0c21; // 0x2556
	13'h12ac: q3 = 16'hca1f; // 0x2558
	13'h12ad: q3 = 16'h808a; // 0x255a
	13'h12ae: q3 = 16'hfd67; // 0x255c
	13'h12af: q3 = 16'h9720; // 0x255e
	13'h12b0: q3 = 16'h30be; // 0x2560
	13'h12b1: q3 = 16'h99ee; // 0x2562
	13'h12b2: q3 = 16'h9650; // 0x2564
	13'h12b3: q3 = 16'h30bf; // 0x2566
	13'h12b4: q3 = 16'h5c80; // 0x2568
	13'h12b5: q3 = 16'hce5b; // 0x256a
	13'h12b6: q3 = 16'h258f; // 0x256c
	13'h12b7: q3 = 16'h4a6f; // 0x256e
	13'h12b8: q3 = 16'hbae9; // 0x2570
	13'h12b9: q3 = 16'h72f8; // 0x2572
	13'h12ba: q3 = 16'hf8d6; // 0x2574
	13'h12bb: q3 = 16'hd033; // 0x2576
	13'h12bc: q3 = 16'hd359; // 0x2578
	13'h12bd: q3 = 16'ha503; // 0x257a
	13'h12be: q3 = 16'had40; // 0x257c
	13'h12bf: q3 = 16'hde19; // 0x257e
	13'h12c0: q3 = 16'h68b2; // 0x2580
	13'h12c1: q3 = 16'h5bbe; // 0x2582
	13'h12c2: q3 = 16'hce5b; // 0x2584
	13'h12c3: q3 = 16'h258e; // 0x2586
	13'h12c4: q3 = 16'h3a6f; // 0x2588
	13'h12c5: q3 = 16'hba1c; // 0x258a
	13'h12c6: q3 = 16'h8096; // 0x258c
	13'h12c7: q3 = 16'hc02e; // 0x258e
	13'h12c8: q3 = 16'ha769; // 0x2590
	13'h12c9: q3 = 16'h6c03; // 0x2592
	13'h12ca: q3 = 16'h902f; // 0x2594
	13'h12cb: q3 = 16'hc32a; // 0x2596
	13'h12cc: q3 = 16'h6da7; // 0x2598
	13'h12cd: q3 = 16'h2f80; // 0x259a
	13'h12ce: q3 = 16'hba9d; // 0x259c
	13'h12cf: q3 = 16'ha587; // 0x259e
	13'h12d0: q3 = 16'h5025; // 0x25a0
	13'h12d1: q3 = 16'hd3e0; // 0x25a2
	13'h12d2: q3 = 16'h86e9; // 0x25a4
	13'h12d3: q3 = 16'h00c3; // 0x25a6
	13'h12d4: q3 = 16'h5ce8; // 0x25a8
	13'h12d5: q3 = 16'h034a; // 0x25aa
	13'h12d6: q3 = 16'h32bf; // 0x25ac
	13'h12d7: q3 = 16'h7034; // 0x25ae
	13'h12d8: q3 = 16'hbc0c; // 0x25b0
	13'h12d9: q3 = 16'hf487; // 0x25b2
	13'h12da: q3 = 16'h2d3e; // 0x25b4
	13'h12db: q3 = 16'hd6e9; // 0x25b6
	13'h12dc: q3 = 16'h00df; // 0x25b8
	13'h12dd: q3 = 16'h5ca6; // 0x25ba
	13'h12de: q3 = 16'h03ad; // 0x25bc
	13'h12df: q3 = 16'h6d03; // 0x25be
	13'h12e0: q3 = 16'h3d21; // 0x25c0
	13'h12e1: q3 = 16'hcb40; // 0x25c2
	13'h12e2: q3 = 16'h24cb; // 0x25c4
	13'h12e3: q3 = 16'h5963; // 0x25c6
	13'h12e4: q3 = 16'hae5b; // 0x25c8
	13'h12e5: q3 = 16'hbe96; // 0x25ca
	13'h12e6: q3 = 16'hc022; // 0x25cc
	13'h12e7: q3 = 16'hbf4b; // 0x25ce
	13'h12e8: q3 = 16'hee02; // 0x25d0
	13'h12e9: q3 = 16'h4940; // 0x25d2
	13'h12ea: q3 = 16'h8efb; // 0x25d4
	13'h12eb: q3 = 16'h6996; // 0x25d6
	13'h12ec: q3 = 16'heeaf; // 0x25d8
	13'h12ed: q3 = 16'h0249; // 0x25da
	13'h12ee: q3 = 16'h40ab; // 0x25dc
	13'h12ef: q3 = 16'h5967; // 0x25de
	13'h12f0: q3 = 16'hbfe0; // 0x25e0
	13'h12f1: q3 = 16'hc2fd; // 0x25e2
	13'h12f2: q3 = 16'h73ce; // 0x25e4
	13'h12f3: q3 = 16'h5e80; // 0x25e6
	13'h12f4: q3 = 16'h8afd; // 0x25e8
	13'h12f5: q3 = 16'h74be; // 0x25ea
	13'h12f6: q3 = 16'he030; // 0x25ec
	13'h12f7: q3 = 16'hbf5c; // 0x25ee
	13'h12f8: q3 = 16'h808e; // 0x25f0
	13'h12f9: q3 = 16'hfb6d; // 0x25f2
	13'h12fa: q3 = 16'h96e8; // 0x25f4
	13'h12fb: q3 = 16'he5cb; // 0x25f6
	13'h12fc: q3 = 16'he0d2; // 0x25f8
	13'h12fd: q3 = 16'h9b65; // 0x25fa
	13'h12fe: q3 = 16'h03e0; // 0x25fc
	13'h12ff: q3 = 16'hea5a; // 0x25fe
	13'h1300: q3 = 16'h7403; // 0x2600
	13'h1301: q3 = 16'he0ce; // 0x2602
	13'h1302: q3 = 16'h59f5; // 0x2604
	13'h1303: q3 = 16'hba4b; // 0x2606
	13'h1304: q3 = 16'hf303; // 0x2608
	13'h1305: q3 = 16'he0d2; // 0x260a
	13'h1306: q3 = 16'h5b70; // 0x260c
	13'h1307: q3 = 16'hcc0f; // 0x260e
	13'h1308: q3 = 16'h8097; // 0x2610
	13'h1309: q3 = 16'h8d32; // 0x2612
	13'h130a: q3 = 16'h8408; // 0x2614
	13'h130b: q3 = 16'he8d6; // 0x2616
	13'h130c: q3 = 16'h3ac0; // 0x2618
	13'h130d: q3 = 16'h8778; // 0x261a
	13'h130e: q3 = 16'h7292; // 0x261c
	13'h130f: q3 = 16'h593e; // 0x261e
	13'h1310: q3 = 16'h978d; // 0x2620
	13'h1311: q3 = 16'h3284; // 0x2622
	13'h1312: q3 = 16'h08e8; // 0x2624
	13'h1313: q3 = 16'hd63a; // 0x2626
	13'h1314: q3 = 16'hc09e; // 0x2628
	13'h1315: q3 = 16'h98b4; // 0x262a
	13'h1316: q3 = 16'h1f3f; // 0x262c
	13'h1317: q3 = 16'h80ce; // 0x262e
	13'h1318: q3 = 16'h5027; // 0x2630
	13'h1319: q3 = 16'h86e8; // 0x2632
	13'h131a: q3 = 16'h40d6; // 0x2634
	13'h131b: q3 = 16'he023; // 0x2636
	13'h131c: q3 = 16'ha358; // 0x2638
	13'h131d: q3 = 16'heb02; // 0x263a
	13'h131e: q3 = 16'h5e34; // 0x263c
	13'h131f: q3 = 16'hca1f; // 0x263e
	13'h1320: q3 = 16'h808e; // 0x2640
	13'h1321: q3 = 16'h8d63; // 0x2642
	13'h1322: q3 = 16'hac0c; // 0x2644
	13'h1323: q3 = 16'hf5c3; // 0x2646
	13'h1324: q3 = 16'h0b25; // 0x2648
	13'h1325: q3 = 16'hb65b; // 0x264a
	13'h1326: q3 = 16'hb486; // 0x264c
	13'h1327: q3 = 16'h9ca5; // 0x264e
	13'h1328: q3 = 16'h0249; // 0x2650
	13'h1329: q3 = 16'h6397; // 0x2652
	13'h132a: q3 = 16'h2ba5; // 0x2654
	13'h132b: q3 = 16'hf887; // 0x2656
	13'h132c: q3 = 16'h403e; // 0x2658
	13'h132d: q3 = 16'h8a5a; // 0x265a
	13'h132e: q3 = 16'h40f8; // 0x265c
	13'h132f: q3 = 16'h840b; // 0x265e
	13'h1330: q3 = 16'h2fcc; // 0x2660
	13'h1331: q3 = 16'h0f80; // 0x2662
	13'h1332: q3 = 16'h840f; // 0x2664
	13'h1333: q3 = 16'h8041; // 0x2666
	13'h1334: q3 = 16'h0030; // 0x2668
	13'h1335: q3 = 16'hbe9b; // 0x266a
	13'h1336: q3 = 16'hb4cf; // 0x266c
	13'h1337: q3 = 16'he041; // 0x266e
	13'h1338: q3 = 16'h0f80; // 0x2670
	13'h1339: q3 = 16'h4100; // 0x2672
	13'h133a: q3 = 16'h30d6; // 0x2674
	13'h133b: q3 = 16'hed2f; // 0x2676
	13'h133c: q3 = 16'hcfe0; // 0x2678
	13'h133d: q3 = 16'h4100; // 0x267a
	13'h133e: q3 = 16'h30be; // 0x267c
	13'h133f: q3 = 16'h9bb4; // 0x267e
	13'h1340: q3 = 16'hcfe0; // 0x2680
	13'h1341: q3 = 16'h021b; // 0x2682
	13'h1342: q3 = 16'ha4f8; // 0x2684
	13'h1343: q3 = 16'h035b; // 0x2686
	13'h1344: q3 = 16'ha4f8; // 0x2688
	13'h1345: q3 = 16'h039f; // 0x268a
	13'h1346: q3 = 16'h8002; // 0x268c
	13'h1347: q3 = 16'h5d3e; // 0x268e
	13'h1348: q3 = 16'h8740; // 0x2690
	13'h1349: q3 = 16'h2586; // 0x2692
	13'h134a: q3 = 16'h3a00; // 0x2694
	13'h134b: q3 = 16'hf88a; // 0x2696
	13'h134c: q3 = 16'h5a40; // 0x2698
	13'h134d: q3 = 16'haa59; // 0x269a
	13'h134e: q3 = 16'h25b8; // 0x269c
	13'h134f: q3 = 16'h0f80; // 0x269e
	13'h1350: q3 = 16'h925c; // 0x26a0
	13'h1351: q3 = 16'hf0d6; // 0x26a2
	13'h1352: q3 = 16'h5cc0; // 0x26a4
	13'h1353: q3 = 16'h9250; // 0x26a6
	13'h1354: q3 = 16'h2386; // 0x26a8
	13'h1355: q3 = 16'h4840; // 0x26aa
	13'h1356: q3 = 16'hf887; // 0x26ac
	13'h1357: q3 = 16'h0ca5; // 0x26ae
	13'h1358: q3 = 16'hcc08; // 0x26b0
	13'h1359: q3 = 16'he887; // 0x26b2
	13'h135a: q3 = 16'h1d65; // 0x26b4
	13'h135b: q3 = 16'h03e0; // 0x26b6
	13'h135c: q3 = 16'h4100; // 0x26b8
	13'h135d: q3 = 16'h30be; // 0x26ba
	13'h135e: q3 = 16'h9bb4; // 0x26bc
	13'h135f: q3 = 16'hcfe0; // 0x26be
	13'h1360: q3 = 16'h410f; // 0x26c0
	13'h1361: q3 = 16'h8041; // 0x26c2
	13'h1362: q3 = 16'h0030; // 0x26c4
	13'h1363: q3 = 16'hd6ed; // 0x26c6
	13'h1364: q3 = 16'h2fcf; // 0x26c8
	13'h1365: q3 = 16'he041; // 0x26ca
	13'h1366: q3 = 16'h0f80; // 0x26cc
	13'h1367: q3 = 16'h021b; // 0x26ce
	13'h1368: q3 = 16'ha4f8; // 0x26d0
	13'h1369: q3 = 16'h035b; // 0x26d2
	13'h136a: q3 = 16'ha4f8; // 0x26d4
	13'h136b: q3 = 16'h039f; // 0x26d6
	13'h136c: q3 = 16'h8002; // 0x26d8
	13'h136d: q3 = 16'h5d00; // 0x26da
	13'h136e: q3 = 16'hc2fd; // 0x26dc
	13'h136f: q3 = 16'h72f8; // 0x26de
	13'h1370: q3 = 16'h9afc; // 0x26e0
	13'h1371: q3 = 16'h80cf; // 0x26e2
	13'h1372: q3 = 16'h4872; // 0x26e4
	13'h1373: q3 = 16'hd29b; // 0x26e6
	13'h1374: q3 = 16'ha702; // 0x26e8
	13'h1375: q3 = 16'h1d00; // 0x26ea
	13'h1376: q3 = 16'ha299; // 0x26ec
	13'h1377: q3 = 16'he802; // 0x26ee
	13'h1378: q3 = 16'hc976; // 0x26f0
	13'h1379: q3 = 16'h96cc; // 0x26f2
	13'h137a: q3 = 16'hfe9b; // 0x26f4
	13'h137b: q3 = 16'h5972; // 0x26f6
	13'h137c: q3 = 16'h033d; // 0x26f8
	13'h137d: q3 = 16'h21cb; // 0x26fa
	13'h137e: q3 = 16'h4022; // 0x26fc
	13'h137f: q3 = 16'h9690; // 0x26fe
	13'h1380: q3 = 16'h28be; // 0x2700
	13'h1381: q3 = 16'h896e; // 0x2702
	13'h1382: q3 = 16'h033d; // 0x2704
	13'h1383: q3 = 16'h359a; // 0x2706
	13'h1384: q3 = 16'h5bbe; // 0x2708
	13'h1385: q3 = 16'h86c0; // 0x270a
	13'h1386: q3 = 16'h23be; // 0x270c
	13'h1387: q3 = 16'hd96e; // 0x270e
	13'h1388: q3 = 16'hea1c; // 0x2710
	13'h1389: q3 = 16'h8084; // 0x2712
	13'h138a: q3 = 16'h086c; // 0x2714
	13'h138b: q3 = 16'hd2fc; // 0x2716
	13'h138c: q3 = 16'hc0ba; // 0x2718
	13'h138d: q3 = 16'h9da5; // 0x271a
	13'h138e: q3 = 16'hb25c; // 0x271c
	13'h138f: q3 = 16'hfe8e; // 0x271e
	13'h1390: q3 = 16'hfb6d; // 0x2720
	13'h1391: q3 = 16'h96e8; // 0x2722
	13'h1392: q3 = 16'he5c8; // 0x2724
	13'h1393: q3 = 16'h0875; // 0x2726
	13'h1394: q3 = 16'he00b; // 0x2728
	13'h1395: q3 = 16'ha9da; // 0x272a
	13'h1396: q3 = 16'h5875; // 0x272c
	13'h1397: q3 = 16'he009; // 0x272e
	13'h1398: q3 = 16'h6c97; // 0x2730
	13'h1399: q3 = 16'h6973; // 0x2732
	13'h139a: q3 = 16'hf8a6; // 0x2734
	13'h139b: q3 = 16'hed32; // 0x2736
	13'h139c: q3 = 16'hbe4d; // 0x2738
	13'h139d: q3 = 16'h63a6; // 0x273a
	13'h139e: q3 = 16'he9ce; // 0x273c
	13'h139f: q3 = 16'h38ef; // 0x273e
	13'h13a0: q3 = 16'h80de; // 0x2740
	13'h13a1: q3 = 16'h9c80; // 0x2742
	13'h13a2: q3 = 16'hcf49; // 0x2744
	13'h13a3: q3 = 16'h6cb2; // 0x2746
	13'h13a4: q3 = 16'h5b80; // 0x2748
	13'h13a5: q3 = 16'hdafc; // 0x274a
	13'h13a6: q3 = 16'h8e38; // 0x274c
	13'h13a7: q3 = 16'hef80; // 0x274e
	13'h13a8: q3 = 16'hc329; // 0x2750
	13'h13a9: q3 = 16'h7396; // 0x2752
	13'h13aa: q3 = 16'hed21; // 0x2754
	13'h13ab: q3 = 16'hb6fc; // 0x2756
	13'h13ac: q3 = 16'hce38; // 0x2758
	13'h13ad: q3 = 16'hef80; // 0x275a
	13'h13ae: q3 = 16'hc329; // 0x275c
	13'h13af: q3 = 16'h7396; // 0x275e
	13'h13b0: q3 = 16'hed21; // 0x2760
	13'h13b1: q3 = 16'hbb43; // 0x2762
	13'h13b2: q3 = 16'h8e3b; // 0x2764
	13'h13b3: q3 = 16'he0cf; // 0x2766
	13'h13b4: q3 = 16'h4872; // 0x2768
	13'h13b5: q3 = 16'hca9b; // 0x276a
	13'h13b6: q3 = 16'ha738; // 0x276c
	13'h13b7: q3 = 16'he3be; // 0x276e
	13'h13b8: q3 = 16'ha6e0; // 0x2770
	13'h13b9: q3 = 16'h2497; // 0x2772
	13'h13ba: q3 = 16'h2028; // 0x2774
	13'h13bb: q3 = 16'h875c; // 0x2776
	13'h13bc: q3 = 16'h34ca; // 0x2778
	13'h13bd: q3 = 16'hfb2c; // 0x277a
	13'h13be: q3 = 16'h94e3; // 0x277c
	13'h13bf: q3 = 16'h8ef8; // 0x277e
	13'h13c0: q3 = 16'h96c0; // 0x2780
	13'h13c1: q3 = 16'h30ca; // 0x2782
	13'h13c2: q3 = 16'hfd21; // 0x2784
	13'h13c3: q3 = 16'h9efb; // 0x2786
	13'h13c4: q3 = 16'ha9cf; // 0x2788
	13'h13c5: q3 = 16'h484e; // 0x278a
	13'h13c6: q3 = 16'h38ef; // 0x278c
	13'h13c7: q3 = 16'h809a; // 0x278e
	13'h13c8: q3 = 16'h99f5; // 0x2790
	13'h13c9: q3 = 16'hca1b; // 0x2792
	13'h13ca: q3 = 16'hb438; // 0x2794
	13'h13cb: q3 = 16'he3be; // 0x2796
	13'h13cc: q3 = 16'hcf48; // 0x2798
	13'h13cd: q3 = 16'h7902; // 0x279a
	13'h13ce: q3 = 16'h1de1; // 0x279c
	13'h13cf: q3 = 16'he409; // 0x279e
	13'h13d0: q3 = 16'hb2be; // 0x27a0
	13'h13d1: q3 = 16'hd023; // 0x27a2
	13'h13d2: q3 = 16'ha259; // 0x27a4
	13'h13d3: q3 = 16'hb3f8; // 0x27a6
	13'h13d4: q3 = 16'h8e89; // 0x27a8
	13'h13d5: q3 = 16'h66ae; // 0x27aa
	13'h13d6: q3 = 16'hf963; // 0x27ac
	13'h13d7: q3 = 16'ha250; // 0x27ae
	13'h13d8: q3 = 16'h2d96; // 0x27b0
	13'h13d9: q3 = 16'h9925; // 0x27b2
	13'h13da: q3 = 16'hbbe0; // 0x27b4
	13'h13db: q3 = 16'hb61b; // 0x27b6
	13'h13dc: q3 = 16'hb496; // 0x27b8
	13'h13dd: q3 = 16'he9e1; // 0x27ba
	13'h13de: q3 = 16'hce50; // 0x27bc
	13'h13df: q3 = 16'h21b2; // 0x27be
	13'h13e0: q3 = 16'h5aa1; // 0x27c0
	13'h13e1: q3 = 16'h92f0; // 0x27c2
	13'h13e2: q3 = 16'h2494; // 0x27c4
	13'h13e3: q3 = 16'h0b2f; // 0x27c6
	13'h13e4: q3 = 16'hcc08; // 0x27c8
	13'h13e5: q3 = 16'he896; // 0x27ca
	13'h13e6: q3 = 16'h6cfe; // 0x27cc
	13'h13e7: q3 = 16'hca5c; // 0x27ce
	13'h13e8: q3 = 16'hf497; // 0x27d0
	13'h13e9: q3 = 16'ha02c; // 0x27d2
	13'h13ea: q3 = 16'hbe9b; // 0x27d4
	13'h13eb: q3 = 16'h8092; // 0x27d6
	13'h13ec: q3 = 16'h5cc0; // 0x27d8
	13'h13ed: q3 = 16'h8e89; // 0x27da
	13'h13ee: q3 = 16'h66cf; // 0x27dc
	13'h13ef: q3 = 16'he0f8; // 0x27de
	13'h13f0: q3 = 16'hf88e; // 0x27e0
	13'h13f1: q3 = 16'hfb61; // 0x27e2
	13'h13f2: q3 = 16'hce50; // 0x27e4
	13'h13f3: q3 = 16'h25b0; // 0x27e6
	13'h13f4: q3 = 16'h0a25; // 0x27e8
	13'h13f5: q3 = 16'hb219; // 0x27ea
	13'h13f6: q3 = 16'h2ff8; // 0x27ec
	13'h13f7: q3 = 16'hb61b; // 0x27ee
	13'h13f8: q3 = 16'ha797; // 0x27f0
	13'h13f9: q3 = 16'ha02c; // 0x27f2
	13'h13fa: q3 = 16'h8409; // 0x27f4
	13'h13fb: q3 = 16'hec86; // 0x27f6
	13'h13fc: q3 = 16'h397e; // 0x27f8
	13'h13fd: q3 = 16'h961d; // 0x27fa
	13'h13fe: q3 = 16'h00d2; // 0x27fc
	13'h13ff: q3 = 16'h8940; // 0x27fe
	13'h1400: q3 = 16'h8efb; // 0x2800
	13'h1401: q3 = 16'ha502; // 0x2802
	13'h1402: q3 = 16'h2966; // 0x2804
	13'h1403: q3 = 16'hbf29; // 0x2806
	13'h1404: q3 = 16'h40a7; // 0x2808
	13'h1405: q3 = 16'h402d; // 0x280a
	13'h1406: q3 = 16'h96cd; // 0x280c
	13'h1407: q3 = 16'h33f8; // 0x280e
	13'h1408: q3 = 16'hde19; // 0x2810
	13'h1409: q3 = 16'ha696; // 0x2812
	13'h140a: q3 = 16'hc036; // 0x2814
	13'h140b: q3 = 16'hbf2b; // 0x2816
	13'h140c: q3 = 16'h40ce; // 0x2818
	13'h140d: q3 = 16'h3a2d; // 0x281a
	13'h140e: q3 = 16'h96ce; // 0x281c
	13'h140f: q3 = 16'ha5b8; // 0x281e
	13'h1410: q3 = 16'h0973; // 0x2820
	13'h1411: q3 = 16'hce5b; // 0x2822
	13'h1412: q3 = 16'hbe86; // 0x2824
	13'h1413: q3 = 16'hed25; // 0x2826
	13'h1414: q3 = 16'hcc09; // 0x2828
	13'h1415: q3 = 16'h2503; // 0x282a
	13'h1416: q3 = 16'h1d65; // 0x282c
	13'h1417: q3 = 16'h0339; // 0x282e
	13'h1418: q3 = 16'h409b; // 0x2830
	13'h1419: q3 = 16'h5ba4; // 0x2832
	13'h141a: q3 = 16'h87e0; // 0x2834
	13'h141b: q3 = 16'h8768; // 0x2836
	13'h141c: q3 = 16'h6ed0; // 0x2838
	13'h141d: q3 = 16'h0c75; // 0x283a
	13'h141e: q3 = 16'h1e5b; // 0x283c
	13'h141f: q3 = 16'h2c94; // 0x283e
	13'h1420: q3 = 16'h09af; // 0x2840
	13'h1421: q3 = 16'hba49; // 0x2842
	13'h1422: q3 = 16'h7ec2; // 0x2844
	13'h1423: q3 = 16'hfa6e; // 0x2846
	13'h1424: q3 = 16'hd336; // 0x2848
	13'h1425: q3 = 16'h8001; // 0x284a
	13'h1426: q3 = 16'h5410; // 0x284c
	13'h1427: q3 = 16'h2ac9; // 0x284e
	13'h1428: q3 = 16'h7696; // 0x2850
	13'h1429: q3 = 16'hcf80; // 0x2852
	13'h142a: q3 = 16'hc35b; // 0x2854
	13'h142b: q3 = 16'habd2; // 0x2856
	13'h142c: q3 = 16'h5680; // 0x2858
	13'h142d: q3 = 16'h0154; // 0x285a
	13'h142e: q3 = 16'h102b; // 0x285c
	13'h142f: q3 = 16'h3d35; // 0x285e
	13'h1430: q3 = 16'h9a5f; // 0x2860
	13'h1431: q3 = 16'h80c3; // 0x2862
	13'h1432: q3 = 16'h5bb4; // 0x2864
	13'h1433: q3 = 16'hbf36; // 0x2866
	13'h1434: q3 = 16'h8001; // 0x2868
	13'h1435: q3 = 16'h5410; // 0x286a
	13'h1436: q3 = 16'h00a0; // 0x286c
	13'h1437: q3 = 16'h2ed6; // 0x286e
	13'h1438: q3 = 16'hd972; // 0x2870
	13'h1439: q3 = 16'hbc09; // 0x2872
	13'h143a: q3 = 16'h2502; // 0x2874
	13'h143b: q3 = 16'hea76; // 0x2876
	13'h143c: q3 = 16'h96cf; // 0x2878
	13'h143d: q3 = 16'h80c2; // 0x287a
	13'h143e: q3 = 16'hfa6e; // 0x287c
	13'h143f: q3 = 16'hd336; // 0x287e
	13'h1440: q3 = 16'h8001; // 0x2880
	13'h1441: q3 = 16'h5410; // 0x2882
	13'h1442: q3 = 16'h2aea; // 0x2884
	13'h1443: q3 = 16'h7696; // 0x2886
	13'h1444: q3 = 16'h1d7e; // 0x2888
	13'h1445: q3 = 16'hc2cd; // 0x288a
	13'h1446: q3 = 16'h7301; // 0x288c
	13'h1447: q3 = 16'h1410; // 0x288e
	13'h1448: q3 = 16'h026b; // 0x2890
	13'h1449: q3 = 16'hf202; // 0x2892
	13'h144a: q3 = 16'h5863; // 0x2894
	13'h144b: q3 = 16'ha009; // 0x2896
	13'h144c: q3 = 16'hafbe; // 0x2898
	13'h144d: q3 = 16'h4f80; // 0x289a
	13'h144e: q3 = 16'hc2cd; // 0x289c
	13'h144f: q3 = 16'h7301; // 0x289e
	13'h1450: q3 = 16'h1410; // 0x28a0
	13'h1451: q3 = 16'h026d; // 0x28a2
	13'h1452: q3 = 16'h65c8; // 0x28a4
	13'h1453: q3 = 16'h0aa5; // 0x28a6
	13'h1454: q3 = 16'h925c; // 0x28a8
	13'h1455: q3 = 16'hc097; // 0x28aa
	13'h1456: q3 = 16'h3ce5; // 0x28ac
	13'h1457: q3 = 16'hbbe0; // 0x28ae
	13'h1458: q3 = 16'hb61c; // 0x28b0
	13'h1459: q3 = 16'hc045; // 0x28b2
	13'h145a: q3 = 16'h0400; // 0x28b4
	13'h145b: q3 = 16'hc35b; // 0x28b6
	13'h145c: q3 = 16'hb4bf; // 0x28b8
	13'h145d: q3 = 16'h3030; // 0x28ba
	13'h145e: q3 = 16'hbf20; // 0x28bc
	13'h145f: q3 = 16'h2386; // 0x28be
	13'h1460: q3 = 16'h4840; // 0x28c0
	13'h1461: q3 = 16'h86ca; // 0x28c2
	13'h1462: q3 = 16'h6d96; // 0x28c4
	13'h1463: q3 = 16'hed2f; // 0x28c6
	13'h1464: q3 = 16'hf8c2; // 0x28c8
	13'h1465: q3 = 16'hcd73; // 0x28ca
	13'h1466: q3 = 16'h0114; // 0x28cc
	13'h1467: q3 = 16'h1003; // 0x28ce
	13'h1468: q3 = 16'h0bf5; // 0x28d0
	13'h1469: q3 = 16'hc808; // 0x28d2
	13'h146a: q3 = 16'he887; // 0x28d4
	13'h146b: q3 = 16'h1d65; // 0x28d6
	13'h146c: q3 = 16'h021b; // 0x28d8
	13'h146d: q3 = 16'h29b6; // 0x28da
	13'h146e: q3 = 16'h5bb4; // 0x28dc
	13'h146f: q3 = 16'hf8f8; // 0x28de
	13'h1470: q3 = 16'hf8ce; // 0x28e0
	13'h1471: q3 = 16'h5027; // 0x28e2
	13'h1472: q3 = 16'h86e8; // 0x28e4
	13'h1473: q3 = 16'h4045; // 0x28e6
	13'h1474: q3 = 16'h040d; // 0x28e8
	13'h1475: q3 = 16'h4504; // 0x28ea
	13'h1476: q3 = 16'h1003; // 0x28ec
	13'h1477: q3 = 16'h0d6e; // 0x28ee
	13'h1478: q3 = 16'hd2fc; // 0x28f0
	13'h1479: q3 = 16'hfef8; // 0x28f2
	13'h147a: q3 = 16'ha29d; // 0x28f4
	13'h147b: q3 = 16'h008e; // 0x28f6
	13'h147c: q3 = 16'h8966; // 0x28f8
	13'h147d: q3 = 16'hcc0d; // 0x28fa
	13'h147e: q3 = 16'he9d2; // 0x28fc
	13'h147f: q3 = 16'h8026; // 0x28fe
	13'h1480: q3 = 16'hbef9; // 0x2900
	13'h1481: q3 = 16'h3e8e; // 0x2902
	13'h1482: q3 = 16'h8966; // 0x2904
	13'h1483: q3 = 16'hcc0b; // 0x2906
	13'h1484: q3 = 16'h69d0; // 0x2908
	13'h1485: q3 = 16'h0973; // 0x290a
	13'h1486: q3 = 16'hce5b; // 0x290c
	13'h1487: q3 = 16'h80d3; // 0x290e
	13'h1488: q3 = 16'h2966; // 0x2910
	13'h1489: q3 = 16'h9a5b; // 0x2912
	13'h148a: q3 = 16'hbe8e; // 0x2914
	13'h148b: q3 = 16'h1921; // 0x2916
	13'h148c: q3 = 16'h0369; // 0x2918
	13'h148d: q3 = 16'h7a03; // 0x291a
	13'h148e: q3 = 16'h1d65; // 0x291c
	13'h148f: q3 = 16'h0339; // 0x291e
	13'h1490: q3 = 16'h4086; // 0x2920
	13'h1491: q3 = 16'h3a65; // 0x2922
	13'h1492: q3 = 16'hcb48; // 0x2924
	13'h1493: q3 = 16'h7e45; // 0x2926
	13'h1494: q3 = 16'h040d; // 0x2928
	13'h1495: q3 = 16'h4504; // 0x292a
	13'h1496: q3 = 16'h1003; // 0x292c
	13'h1497: q3 = 16'h0be9; // 0x292e
	13'h1498: q3 = 16'hbb4c; // 0x2930
	13'h1499: q3 = 16'hc08e; // 0x2932
	13'h149a: q3 = 16'h8871; // 0x2934
	13'h149b: q3 = 16'hd650; // 0x2936
	13'h149c: q3 = 16'h26be; // 0x2938
	13'h149d: q3 = 16'h9cc0; // 0x293a
	13'h149e: q3 = 16'hc759; // 0x293c
	13'h149f: q3 = 16'h7e45; // 0x293e
	13'h14a0: q3 = 16'h040d; // 0x2940
	13'h14a1: q3 = 16'h4504; // 0x2942
	13'h14a2: q3 = 16'h1003; // 0x2944
	13'h14a3: q3 = 16'h0be9; // 0x2946
	13'h14a4: q3 = 16'hbb4c; // 0x2948
	13'h14a5: q3 = 16'hfe45; // 0x294a
	13'h14a6: q3 = 16'h040d; // 0x294c
	13'h14a7: q3 = 16'h4504; // 0x294e
	13'h14a8: q3 = 16'h1003; // 0x2950
	13'h14a9: q3 = 16'h0d6e; // 0x2952
	13'h14aa: q3 = 16'haf49; // 0x2954
	13'h14ab: q3 = 16'h7e84; // 0x2956
	13'h14ac: q3 = 16'h0b2f; // 0x2958
	13'h14ad: q3 = 16'hcc08; // 0x295a
	13'h14ae: q3 = 16'he896; // 0x295c
	13'h14af: q3 = 16'h6cc0; // 0x295e
	13'h14b0: q3 = 16'h8efb; // 0x2960
	13'h14b1: q3 = 16'h8086; // 0x2962
	13'h14b2: q3 = 16'hca6d; // 0x2964
	13'h14b3: q3 = 16'h96ed; // 0x2966
	13'h14b4: q3 = 16'h2fcf; // 0x2968
	13'h14b5: q3 = 16'he0da; // 0x296a
	13'h14b6: q3 = 16'hfd73; // 0x296c
	13'h14b7: q3 = 16'h026c; // 0x296e
	13'h14b8: q3 = 16'ha1c3; // 0x2970
	13'h14b9: q3 = 16'h097a; // 0x2972
	13'h14ba: q3 = 16'h023a; // 0x2974
	13'h14bb: q3 = 16'h259b; // 0x2976
	13'h14bc: q3 = 16'h3021; // 0x2978
	13'h14bd: q3 = 16'hda58; // 0x297a
	13'h14be: q3 = 16'hc086; // 0x297c
	13'h14bf: q3 = 16'hca6d; // 0x297e
	13'h14c0: q3 = 16'h96ed; // 0x2980
	13'h14c1: q3 = 16'h3e87; // 0x2982
	13'h14c2: q3 = 16'h2b40; // 0x2984
	13'h14c3: q3 = 16'hc2fa; // 0x2986
	13'h14c4: q3 = 16'h6ed3; // 0x2988
	13'h14c5: q3 = 16'h3029; // 0x298a
	13'h14c6: q3 = 16'hb809; // 0x298c
	13'h14c7: q3 = 16'h29ca; // 0x298e
	13'h14c8: q3 = 16'h58f4; // 0x2990
	13'h14c9: q3 = 16'ha6fb; // 0x2992
	13'h14ca: q3 = 16'hbe87; // 0x2994
	13'h14cb: q3 = 16'h2b40; // 0x2996
	13'h14cc: q3 = 16'hea5a; // 0x2998
	13'h14cd: q3 = 16'h67d3; // 0x299a
	13'h14ce: q3 = 16'he096; // 0x299c
	13'h14cf: q3 = 16'hc022; // 0x299e
	13'h14d0: q3 = 16'hca1e; // 0x29a0
	13'h14d1: q3 = 16'haf02; // 0x29a2
	13'h14d2: q3 = 16'h1c35; // 0x29a4
	13'h14d3: q3 = 16'hbb48; // 0x29a6
	13'h14d4: q3 = 16'h4096; // 0x29a8
	13'h14d5: q3 = 16'he025; // 0x29aa
	13'h14d6: q3 = 16'hb00c; // 0x29ac
	13'h14d7: q3 = 16'he5bb; // 0x29ae
	13'h14d8: q3 = 16'h4a64; // 0x29b0
	13'h14d9: q3 = 16'hbc09; // 0x29b2
	13'h14da: q3 = 16'h6ef8; // 0x29b4
	13'h14db: q3 = 16'h8b28; // 0x29b6
	13'h14dc: q3 = 16'h7303; // 0x29b8
	13'h14dd: q3 = 16'h0be9; // 0x29ba
	13'h14de: q3 = 16'hbb49; // 0x29bc
	13'h14df: q3 = 16'h4096; // 0x29be
	13'h14e0: q3 = 16'he024; // 0x29c0
	13'h14e1: q3 = 16'ha729; // 0x29c2
	13'h14e2: q3 = 16'h63d2; // 0x29c4
	13'h14e3: q3 = 16'h9bee; // 0x29c6
	13'h14e4: q3 = 16'hf8be; // 0x29c8
	13'h14e5: q3 = 16'h6034; // 0x29ca
	13'h14e6: q3 = 16'ha32b; // 0x29cc
	13'h14e7: q3 = 16'hf7f8; // 0x29ce
	13'h14e8: q3 = 16'ha6e0; // 0x29d0
	13'h14e9: q3 = 16'h37d7; // 0x29d2
	13'h14ea: q3 = 16'h29b2; // 0x29d4
	13'h14eb: q3 = 16'ha63a; // 0x29d6
	13'h14ec: q3 = 16'h34d6; // 0x29d8
	13'h14ed: q3 = 16'he9fe; // 0x29da
	13'h14ee: q3 = 16'hc759; // 0x29dc
	13'h14ef: q3 = 16'h40ce; // 0x29de
	13'h14f0: q3 = 16'h502c; // 0x29e0
	13'h14f1: q3 = 16'h86ee; // 0x29e2
	13'h14f2: q3 = 16'ha102; // 0x29e4
	13'h14f3: q3 = 16'h5b00; // 0x29e6
	13'h14f4: q3 = 16'h86ca; // 0x29e8
	13'h14f5: q3 = 16'h6d96; // 0x29ea
	13'h14f6: q3 = 16'hed2f; // 0x29ec
	13'h14f7: q3 = 16'hf893; // 0x29ee
	13'h14f8: q3 = 16'h502c; // 0x29f0
	13'h14f9: q3 = 16'h86e8; // 0x29f2
	13'h14fa: q3 = 16'he5f8; // 0x29f4
	13'h14fb: q3 = 16'h876b; // 0x29f6
	13'h14fc: q3 = 16'he990; // 0x29f8
	13'h14fd: q3 = 16'h09af; // 0x29fa
	13'h14fe: q3 = 16'hbe40; // 0x29fc
	13'h14ff: q3 = 16'h34a3; // 0x29fe
	13'h1500: q3 = 16'h2bf7; // 0x2a00
	13'h1501: q3 = 16'hb808; // 0x2a02
	13'h1502: q3 = 16'hb902; // 0x2a04
	13'h1503: q3 = 16'h3a25; // 0x2a06
	13'h1504: q3 = 16'h9b3f; // 0x2a08
	13'h1505: q3 = 16'h80da; // 0x2a0a
	13'h1506: q3 = 16'hfb80; // 0x2a0c
	13'h1507: q3 = 16'h8e89; // 0x2a0e
	13'h1508: q3 = 16'h66cc; // 0x2a10
	13'h1509: q3 = 16'h09e5; // 0x2a12
	13'h150a: q3 = 16'hdefc; // 0x2a14
	13'h150b: q3 = 16'ha696; // 0x2a16
	13'h150c: q3 = 16'he973; // 0x2a18
	13'h150d: q3 = 16'hf897; // 0x2a1a
	13'h150e: q3 = 16'h3c75; // 0x2a1c
	13'h150f: q3 = 16'ha769; // 0x2a1e
	13'h1510: q3 = 16'h4096; // 0x2a20
	13'h1511: q3 = 16'hc021; // 0x2a22
	13'h1512: q3 = 16'hb29b; // 0x2a24
	13'h1513: q3 = 16'h65bb; // 0x2a26
	13'h1514: q3 = 16'h4bfe; // 0x2a28
	13'h1515: q3 = 16'h976a; // 0x2a2a
	13'h1516: q3 = 16'h7497; // 0x2a2c
	13'h1517: q3 = 16'ha021; // 0x2a2e
	13'h1518: q3 = 16'hb29b; // 0x2a30
	13'h1519: q3 = 16'h65bb; // 0x2a32
	13'h151a: q3 = 16'h4cfe; // 0x2a34
	13'h151b: q3 = 16'hf897; // 0x2a36
	13'h151c: q3 = 16'h3ce5; // 0x2a38
	13'h151d: q3 = 16'hb80d; // 0x2a3a
	13'h151e: q3 = 16'ha5ca; // 0x2a3c
	13'h151f: q3 = 16'hd969; // 0x2a3e
	13'h1520: q3 = 16'h925b; // 0x2a40
	13'h1521: q3 = 16'hbeb2; // 0x2a42
	13'h1522: q3 = 16'h1bba; // 0x2a44
	13'h1523: q3 = 16'h864b; // 0x2a46
	13'h1524: q3 = 16'hc0c2; // 0x2a48
	13'h1525: q3 = 16'hfc80; // 0x2a4a
	13'h1526: q3 = 16'hb2fc; // 0x2a4c
	13'h1527: q3 = 16'hc08e; // 0x2a4e
	13'h1528: q3 = 16'h8966; // 0x2a50
	13'h1529: q3 = 16'hcfe0; // 0x2a52
	13'h152a: q3 = 16'hb21b; // 0x2a54
	13'h152b: q3 = 16'ha397; // 0x2a56
	13'h152c: q3 = 16'h3030; // 0x2a58
	13'h152d: q3 = 16'h8720; // 0x2a5a
	13'h152e: q3 = 16'h23a2; // 0x2a5c
	13'h152f: q3 = 16'h59b3; // 0x2a5e
	13'h1530: q3 = 16'hf88e; // 0x2a60
	13'h1531: q3 = 16'h8966; // 0x2a62
	13'h1532: q3 = 16'h0268; // 0x2a64
	13'h1533: q3 = 16'h6cb3; // 0x2a66
	13'h1534: q3 = 16'h3029; // 0x2a68
	13'h1535: q3 = 16'hbb4b; // 0x2a6a
	13'h1536: q3 = 16'hc0a2; // 0x2a6c
	13'h1537: q3 = 16'hfb25; // 0x2a6e
	13'h1538: q3 = 16'hf88e; // 0x2a70
	13'h1539: q3 = 16'h8966; // 0x2a72
	13'h153a: q3 = 16'h0268; // 0x2a74
	13'h153b: q3 = 16'h65b2; // 0x2a76
	13'h153c: q3 = 16'hcd00; // 0x2a78
	13'h153d: q3 = 16'ha6ec; // 0x2a7a
	13'h153e: q3 = 16'hc0b2; // 0x2a7c
	13'h153f: q3 = 16'hf8e8; // 0x2a7e
	13'h1540: q3 = 16'hf849; // 0x2a80
	13'h1541: q3 = 16'h0400; // 0x2a82
	13'h1542: q3 = 16'hc35b; // 0x2a84
	13'h1543: q3 = 16'hb4bf; // 0x2a86
	13'h1544: q3 = 16'h3023; // 0x2a88
	13'h1545: q3 = 16'h8648; // 0x2a8a
	13'h1546: q3 = 16'h40da; // 0x2a8c
	13'h1547: q3 = 16'h5e80; // 0x2a8e
	13'h1548: q3 = 16'hc759; // 0x2a90
	13'h1549: q3 = 16'h40d6; // 0x2a92
	13'h154a: q3 = 16'hef80; // 0x2a94
	13'h154b: q3 = 16'h4904; // 0x2a96
	13'h154c: q3 = 16'h00c2; // 0x2a98
	13'h154d: q3 = 16'hfa6e; // 0x2a9a
	13'h154e: q3 = 16'hd330; // 0x2a9c
	13'h154f: q3 = 16'h23a2; // 0x2a9e
	13'h1550: q3 = 16'h1c75; // 0x2aa0
	13'h1551: q3 = 16'h9409; // 0x2aa2
	13'h1552: q3 = 16'hafa7; // 0x2aa4
	13'h1553: q3 = 16'h3031; // 0x2aa6
	13'h1554: q3 = 16'hd47d; // 0x2aa8
	13'h1555: q3 = 16'h6ef8; // 0x2aaa
	13'h1556: q3 = 16'h4904; // 0x2aac
	13'h1557: q3 = 16'h00c2; // 0x2aae
	13'h1558: q3 = 16'hfa6e; // 0x2ab0
	13'h1559: q3 = 16'hd33f; // 0x2ab2
	13'h155a: q3 = 16'h8049; // 0x2ab4
	13'h155b: q3 = 16'h0400; // 0x2ab6
	13'h155c: q3 = 16'hc35b; // 0x2ab8
	13'h155d: q3 = 16'habd2; // 0x2aba
	13'h155e: q3 = 16'h5f80; // 0x2abc
	13'h155f: q3 = 16'h8e89; // 0x2abe
	13'h1560: q3 = 16'h6603; // 0x2ac0
	13'h1561: q3 = 16'h3940; // 0x2ac2
	13'h1562: q3 = 16'h8e19; // 0x2ac4
	13'h1563: q3 = 16'h4092; // 0x2ac6
	13'h1564: q3 = 16'h5bb4; // 0x2ac8
	13'h1565: q3 = 16'hcaf0; // 0x2aca
	13'h1566: q3 = 16'h2494; // 0x2acc
	13'h1567: q3 = 16'h0d6e; // 0x2ace
	13'h1568: q3 = 16'h0219; // 0x2ad0
	13'h1569: q3 = 16'hf5aa; // 0x2ad2
	13'h156a: q3 = 16'h5caf; // 0x2ad4
	13'h156b: q3 = 16'hf88e; // 0x2ad6
	13'h156c: q3 = 16'h8966; // 0x2ad8
	13'h156d: q3 = 16'h025c; // 0x2ada
	13'h156e: q3 = 16'hf403; // 0x2adc
	13'h156f: q3 = 16'h4bed; // 0x2ade
	13'h1570: q3 = 16'h8a50; // 0x2ae0
	13'h1571: q3 = 16'h2486; // 0x2ae2
	13'h1572: q3 = 16'hecc0; // 0x2ae4
	13'h1573: q3 = 16'hd6e0; // 0x2ae6
	13'h1574: q3 = 16'h34ca; // 0x2ae8
	13'h1575: q3 = 16'hfd7e; // 0x2aea
	13'h1576: q3 = 16'hf8f8; // 0x2aec
	13'h1577: q3 = 16'h8f5a; // 0x2aee
	13'h1578: q3 = 16'h6486; // 0x2af0
	13'h1579: q3 = 16'h4bc0; // 0x2af2
	13'h157a: q3 = 16'h8efb; // 0x2af4
	13'h157b: q3 = 16'hbef8; // 0x2af6
	13'h157c: q3 = 16'hde1d; // 0x2af8
	13'h157d: q3 = 16'h23a0; // 0x2afa
	13'h157e: q3 = 16'h0bf5; // 0x2afc
	13'h157f: q3 = 16'hd009; // 0x2afe
	13'h1580: q3 = 16'hafc8; // 0x2b00
	13'h1581: q3 = 16'h0bf0; // 0x2b02
	13'h1582: q3 = 16'h96e0; // 0x2b04
	13'h1583: q3 = 16'h28be; // 0x2b06
	13'h1584: q3 = 16'hc973; // 0x2b08
	13'h1585: q3 = 16'hf886; // 0x2b0a
	13'h1586: q3 = 16'h3a34; // 0x2b0c
	13'h1587: q3 = 16'hd6e9; // 0x2b0e
	13'h1588: q3 = 16'hda00; // 0x2b10
	13'h1589: q3 = 16'h0be6; // 0x2b12
	13'h158a: q3 = 16'h9a5b; // 0x2b14
	13'h158b: q3 = 16'ha502; // 0x2b16
	13'h158c: q3 = 16'hcbe5; // 0x2b18
	13'h158d: q3 = 16'h8e89; // 0x2b1a
	13'h158e: q3 = 16'h72f8; // 0x2b1c
	13'h158f: q3 = 16'hb2fc; // 0x2b1e
	13'h1590: q3 = 16'hc086; // 0x2b20
	13'h1591: q3 = 16'h7d6a; // 0x2b22
	13'h1592: q3 = 16'h972b; // 0x2b24
	13'h1593: q3 = 16'hf302; // 0x2b26
	13'h1594: q3 = 16'h18a9; // 0x2b28
	13'h1595: q3 = 16'h972d; // 0x2b2a
	13'h1596: q3 = 16'h2fcf; // 0x2b2c
	13'h1597: q3 = 16'he087; // 0x2b2e
	13'h1598: q3 = 16'h4d25; // 0x2b30
	13'h1599: q3 = 16'hbb4a; // 0x2b32
	13'h159a: q3 = 16'h6fb8; // 0x2b34
	13'h159b: q3 = 16'h0875; // 0x2b36
	13'h159c: q3 = 16'he00d; // 0x2b38
	13'h159d: q3 = 16'h32bf; // 0x2b3a
	13'h159e: q3 = 16'h5cc0; // 0x2b3c
	13'h159f: q3 = 16'hbf5d; // 0x2b3e
	13'h15a0: q3 = 16'ha5cb; // 0x2b40
	13'h15a1: q3 = 16'h4cfe; // 0x2b42
	13'h15a2: q3 = 16'h4408; // 0x2b44
	13'h15a3: q3 = 16'hf296; // 0x2b46
	13'h15a4: q3 = 16'h4a74; // 0x2b48
	13'h15a5: q3 = 16'hf844; // 0x2b4a
	13'h15a6: q3 = 16'h0cf0; // 0x2b4c
	13'h15a7: q3 = 16'ha65b; // 0x2b4e
	13'h15a8: q3 = 16'h3e44; // 0x2b50
	13'h15a9: q3 = 16'h0ab5; // 0x2b52
	13'h15aa: q3 = 16'h9e19; // 0x2b54
	13'h15ab: q3 = 16'h21f8; // 0x2b56
	13'h15ac: q3 = 16'h4408; // 0x2b58
	13'h15ad: q3 = 16'hf296; // 0x2b5a
	13'h15ae: q3 = 16'h4a74; // 0x2b5c
	13'h15af: q3 = 16'hf802; // 0x2b5e
	13'h15b0: q3 = 16'h3ca5; // 0x2b60
	13'h15b1: q3 = 16'h929d; // 0x2b62
	13'h15b2: q3 = 16'h33f8; // 0x2b64
	13'h15b3: q3 = 16'h033c; // 0x2b66
	13'h15b4: q3 = 16'h2996; // 0x2b68
	13'h15b5: q3 = 16'hc97e; // 0x2b6a
	13'h15b6: q3 = 16'h02ad; // 0x2b6c
	13'h15b7: q3 = 16'h6786; // 0x2b6e
	13'h15b8: q3 = 16'h4873; // 0x2b70
	13'h15b9: q3 = 16'hf802; // 0x2b72
	13'h15ba: q3 = 16'h3ca5; // 0x2b74
	13'h15bb: q3 = 16'h929d; // 0x2b76
	13'h15bc: q3 = 16'h33f8; // 0x2b78
	13'h15bd: q3 = 16'hc329; // 0x2b7a
	13'h15be: q3 = 16'h73cc; // 0x2b7c
	13'h15bf: q3 = 16'h0440; // 0x2b7e
	13'h15c0: q3 = 16'hc2c8; // 0x2b80
	13'h15c1: q3 = 16'h7997; // 0x2b82
	13'h15c2: q3 = 16'h2033; // 0x2b84
	13'h15c3: q3 = 16'hd21c; // 0x2b86
	13'h15c4: q3 = 16'hb4f8; // 0x2b88
	13'h15c5: q3 = 16'h440c; // 0x2b8a
	13'h15c6: q3 = 16'hf0a6; // 0x2b8c
	13'h15c7: q3 = 16'h5b25; // 0x2b8e
	13'h15c8: q3 = 16'hc80c; // 0x2b90
	13'h15c9: q3 = 16'hf487; // 0x2b92
	13'h15ca: q3 = 16'h2d00; // 0x2b94
	13'h15cb: q3 = 16'h932d; // 0x2b96
	13'h15cc: q3 = 16'h658e; // 0x2b98
	13'h15cd: q3 = 16'hb96e; // 0x2b9a
	13'h15ce: q3 = 16'hf8bf; // 0x2b9c
	13'h15cf: q3 = 16'h0ca9; // 0x2b9e
	13'h15d0: q3 = 16'hb69c; // 0x2ba0
	13'h15d1: q3 = 16'h808a; // 0x2ba2
	13'h15d2: q3 = 16'hfd2f; // 0x2ba4
	13'h15d3: q3 = 16'hb80c; // 0x2ba6
	13'h15d4: q3 = 16'h21ca; // 0x2ba8
	13'h15d5: q3 = 16'h1011; // 0x2baa
	13'h15d6: q3 = 16'h02ad; // 0x2bac
	13'h15d7: q3 = 16'h6786; // 0x2bae
	13'h15d8: q3 = 16'h4bf2; // 0x2bb0
	13'h15d9: q3 = 16'hf8c3; // 0x2bb2
	13'h15da: q3 = 16'h2973; // 0x2bb4
	13'h15db: q3 = 16'hce5e; // 0x2bb6
	13'h15dc: q3 = 16'h808a; // 0x2bb8
	13'h15dd: q3 = 16'hfd74; // 0x2bba
	13'h15de: q3 = 16'hbee0; // 0x2bbc
	13'h15df: q3 = 16'h30bf; // 0x2bbe
	13'h15e0: q3 = 16'h5c80; // 0x2bc0
	13'h15e1: q3 = 16'h440a; // 0x2bc2
	13'h15e2: q3 = 16'hafd6; // 0x2bc4
	13'h15e3: q3 = 16'h5d72; // 0x2bc6
	13'h15e4: q3 = 16'hf8c3; // 0x2bc8
	13'h15e5: q3 = 16'h2973; // 0x2bca
	13'h15e6: q3 = 16'hcc04; // 0x2bcc
	13'h15e7: q3 = 16'h40c2; // 0x2bce
	13'h15e8: q3 = 16'hc879; // 0x2bd0
	13'h15e9: q3 = 16'h9720; // 0x2bd2
	13'h15ea: q3 = 16'h2fc8; // 0x2bd4
	13'h15eb: q3 = 16'h0480; // 0x2bd6
	13'h15ec: q3 = 16'hc2c8; // 0x2bd8
	13'h15ed: q3 = 16'h7997; // 0x2bda
	13'h15ee: q3 = 16'h2f80; // 0x2bdc
	13'h15ef: q3 = 16'h440b; // 0x2bde
	13'h15f0: q3 = 16'he497; // 0x2be0
	13'h15f1: q3 = 16'h2012; // 0x2be2
	13'h15f2: q3 = 16'h033c; // 0x2be4
	13'h15f3: q3 = 16'h2996; // 0x2be6
	13'h15f4: q3 = 16'hc972; // 0x2be8
	13'h15f5: q3 = 16'h024c; // 0x2bea
	13'h15f6: q3 = 16'hb596; // 0x2bec
	13'h15f7: q3 = 16'h3ae5; // 0x2bee
	13'h15f8: q3 = 16'hbbe0; // 0x2bf0
	13'h15f9: q3 = 16'hbc04; // 0x2bf2
	13'h15fa: q3 = 16'h80ab; // 0x2bf4
	13'h15fb: q3 = 16'h59e1; // 0x2bf6
	13'h15fc: q3 = 16'h92fc; // 0x2bf8
	13'h15fd: q3 = 16'ha5cf; // 0x2bfa
	13'h15fe: q3 = 16'he0bf; // 0x2bfc
	13'h15ff: q3 = 16'h5012; // 0x2bfe
	13'h1600: q3 = 16'h02ab; // 0x2c00
	13'h1601: q3 = 16'hf597; // 0x2c02
	13'h1602: q3 = 16'h5cb3; // 0x2c04
	13'h1603: q3 = 16'hf8a6; // 0x2c06
	13'h1604: q3 = 16'hece5; // 0x2c08
	13'h1605: q3 = 16'hcb40; // 0x2c0a
	13'h1606: q3 = 16'h23be; // 0x2c0c
	13'h1607: q3 = 16'h9bbe; // 0x2c0e
	13'h1608: q3 = 16'hb759; // 0x2c10
	13'h1609: q3 = 16'h6eea; // 0x2c12
	13'h160a: q3 = 16'h5025; // 0x2c14
	13'h160b: q3 = 16'ha6ed; // 0x2c16
	13'h160c: q3 = 16'he5ca; // 0x2c18
	13'h160d: q3 = 16'h696e; // 0x2c1a
	13'h160e: q3 = 16'hf8a6; // 0x2c1c
	13'h160f: q3 = 16'hece5; // 0x2c1e
	13'h1610: q3 = 16'hcb48; // 0x2c20
	13'h1611: q3 = 16'h7202; // 0x2c22
	13'h1612: q3 = 16'hdbee; // 0x2c24
	13'h1613: q3 = 16'h9648; // 0x2c26
	13'h1614: q3 = 16'h7ea6; // 0x2c28
	13'h1615: q3 = 16'hed32; // 0x2c2a
	13'h1616: q3 = 16'hbe4d; // 0x2c2c
	13'h1617: q3 = 16'h69ce; // 0x2c2e
	13'h1618: q3 = 16'h5e80; // 0x2c30
	13'h1619: q3 = 16'hc299; // 0x2c32
	13'h161a: q3 = 16'h6397; // 0x2c34
	13'h161b: q3 = 16'he09e; // 0x2c36
	13'h161c: q3 = 16'h1b65; // 0x2c38
	13'h161d: q3 = 16'h02fd; // 0x2c3a
	13'h161e: q3 = 16'ha5c8; // 0x2c3c
	13'h161f: q3 = 16'h0c2c; // 0x2c3e
	13'h1620: q3 = 16'h8799; // 0x2c40
	13'h1621: q3 = 16'h7203; // 0x2c42
	13'h1622: q3 = 16'he0cf; // 0x2c44
	13'h1623: q3 = 16'h0a65; // 0x2c46
	13'h1624: q3 = 16'hb009; // 0x2c48
	13'h1625: q3 = 16'hb597; // 0x2c4a
	13'h1626: q3 = 16'h2033; // 0x2c4c
	13'h1627: q3 = 16'hc299; // 0x2c4e
	13'h1628: q3 = 16'h6c97; // 0x2c50
	13'h1629: q3 = 16'h203e; // 0x2c52
	13'h162a: q3 = 16'h9a9b; // 0x2c54
	13'h162b: q3 = 16'h8092; // 0x2c56
	13'h162c: q3 = 16'h502a; // 0x2c58
	13'h162d: q3 = 16'hd659; // 0x2c5a
	13'h162e: q3 = 16'hef03; // 0x2c5c
	13'h162f: q3 = 16'h0872; // 0x2c5e
	13'h1630: q3 = 16'h840a; // 0x2c60
	13'h1631: q3 = 16'hb59e; // 0x2c62
	13'h1632: q3 = 16'h192f; // 0x2c64
	13'h1633: q3 = 16'hc80f; // 0x2c66
	13'h1634: q3 = 16'h80aa; // 0x2c68
	13'h1635: q3 = 16'h5d40; // 0x2c6a
	13'h1636: q3 = 16'hd25c; // 0x2c6c
	13'h1637: q3 = 16'hada6; // 0x2c6e
	13'h1638: q3 = 16'he940; // 0x2c70
	13'h1639: q3 = 16'hc2fd; // 0x2c72
	13'h163a: q3 = 16'h7202; // 0x2c74
	13'h163b: q3 = 16'habf5; // 0x2c76
	13'h163c: q3 = 16'h975c; // 0x2c78
	13'h163d: q3 = 16'h80f8; // 0x2c7a
	13'h163e: q3 = 16'hbf09; // 0x2c7c
	13'h163f: q3 = 16'h6ef8; // 0x2c7e
	13'h1640: q3 = 16'hbe69; // 0x2c80
	13'h1641: q3 = 16'ha5bb; // 0x2c82
	13'h1642: q3 = 16'he086; // 0x2c84
	13'h1643: q3 = 16'h2a65; // 0x2c86
	13'h1644: q3 = 16'hcb4b; // 0x2c88
	13'h1645: q3 = 16'hfebf; // 0x2c8a
	13'h1646: q3 = 16'h5da5; // 0x2c8c
	13'h1647: q3 = 16'hcb4f; // 0x2c8e
	13'h1648: q3 = 16'h808e; // 0x2c90
	13'h1649: q3 = 16'hcbf3; // 0x2c92
	13'h164a: q3 = 16'h964f; // 0x2c94
	13'h164b: q3 = 16'h809e; // 0x2c96
	13'h164c: q3 = 16'h5ce3; // 0x2c98
	13'h164d: q3 = 16'ha2cb; // 0x2c9a
	13'h164e: q3 = 16'hf3ce; // 0x2c9c
	13'h164f: q3 = 16'h5bbe; // 0x2c9e
	13'h1650: q3 = 16'h8e5c; // 0x2ca0
	13'h1651: q3 = 16'hb286; // 0x2ca2
	13'h1652: q3 = 16'h4bfe; // 0x2ca4
	13'h1653: q3 = 16'h9a5c; // 0x2ca6
	13'h1654: q3 = 16'had97; // 0x2ca8
	13'h1655: q3 = 16'he0c3; // 0x2caa
	13'h1656: q3 = 16'h5ce8; // 0x2cac
	13'h1657: q3 = 16'h034a; // 0x2cae
	13'h1658: q3 = 16'h32bf; // 0x2cb0
	13'h1659: q3 = 16'h7034; // 0x2cb2
	13'h165a: q3 = 16'hbc0c; // 0x2cb4
	13'h165b: q3 = 16'he5b2; // 0x2cb6
	13'h165c: q3 = 16'h58f4; // 0x2cb8
	13'h165d: q3 = 16'h02c9; // 0x2cba
	13'h165e: q3 = 16'h74d2; // 0x2cbc
	13'h165f: q3 = 16'h5cbe; // 0x2cbe
	13'h1660: q3 = 16'hdf5c; // 0x2cc0
	13'h1661: q3 = 16'ha602; // 0x2cc2
	13'h1662: q3 = 16'h4cb5; // 0x2cc4
	13'h1663: q3 = 16'h963a; // 0x2cc6
	13'h1664: q3 = 16'he5b9; // 0x2cc8
	13'h1665: q3 = 16'ha000; // 0x2cca
	13'h1666: q3 = 16'h8b58; // 0x2ccc
	13'h1667: q3 = 16'he8cf; // 0x2cce
	13'h1668: q3 = 16'h4862; // 0x2cd0
	13'h1669: q3 = 16'h96ed; // 0x2cd2
	13'h166a: q3 = 16'he1a2; // 0x2cd4
	13'h166b: q3 = 16'hcf80; // 0x2cd6
	13'h166c: q3 = 16'hbf0c; // 0x2cd8
	13'h166d: q3 = 16'ha9b6; // 0x2cda
	13'h166e: q3 = 16'h9c80; // 0x2cdc
	13'h166f: q3 = 16'h8afd; // 0x2cde
	13'h1670: q3 = 16'h2fb8; // 0x2ce0
	13'h1671: q3 = 16'h0c21; // 0x2ce2
	13'h1672: q3 = 16'hca1f; // 0x2ce4
	13'h1673: q3 = 16'h80c2; // 0x2ce6
	13'h1674: q3 = 16'hfd73; // 0x2ce8
	13'h1675: q3 = 16'hce5e; // 0x2cea
	13'h1676: q3 = 16'h808a; // 0x2cec
	13'h1677: q3 = 16'hfd74; // 0x2cee
	13'h1678: q3 = 16'hbee0; // 0x2cf0
	13'h1679: q3 = 16'h30bf; // 0x2cf2
	13'h167a: q3 = 16'h5cbe; // 0x2cf4
	13'h167b: q3 = 16'hf8f8; // 0x2cf6
	13'h167c: q3 = 16'h9738; // 0x2cf8
	13'h167d: q3 = 16'hef9e; // 0x2cfa
	13'h167e: q3 = 16'h5c80; // 0x2cfc
	13'h167f: q3 = 16'hb25d; // 0x2cfe
	13'h1680: q3 = 16'h3287; // 0x2d00
	13'h1681: q3 = 16'h3f80; // 0x2d02
	13'h1682: q3 = 16'hce5b; // 0x2d04
	13'h1683: q3 = 16'h258f; // 0x2d06
	13'h1684: q3 = 16'h4a6f; // 0x2d08
	13'h1685: q3 = 16'hbae9; // 0x2d0a
	13'h1686: q3 = 16'h7202; // 0x2d0c
	13'h1687: q3 = 16'hc974; // 0x2d0e
	13'h1688: q3 = 16'hd329; // 0x2d10
	13'h1689: q3 = 16'h7e9f; // 0x2d12
	13'h168a: q3 = 16'h2961; // 0x2d14
	13'h168b: q3 = 16'hd00c; // 0x2d16
	13'h168c: q3 = 16'he3bf; // 0x2d18
	13'h168d: q3 = 16'h2940; // 0x2d1a
	13'h168e: q3 = 16'hc2c8; // 0x2d1c
	13'h168f: q3 = 16'h7997; // 0x2d1e
	13'h1690: q3 = 16'h203e; // 0x2d20
	13'h1691: q3 = 16'hd2fb; // 0x2d22
	13'h1692: q3 = 16'h2c94; // 0x2d24
	13'h1693: q3 = 16'h0c35; // 0x2d26
	13'h1694: q3 = 16'hbabd; // 0x2d28
	13'h1695: q3 = 16'h25ea; // 0x2d2a
	13'h1696: q3 = 16'h1a2c; // 0x2d2c
	13'h1697: q3 = 16'h300b; // 0x2d2e
	13'h1698: q3 = 16'hb23b; // 0x2d30
	13'h1699: q3 = 16'he012; // 0x2d32
	13'h169a: q3 = 16'h5e23; // 0x2d34
	13'h169b: q3 = 16'h96c9; // 0x2d36
	13'h169c: q3 = 16'h6ed2; // 0x2d38
	13'h169d: q3 = 16'h5030; // 0x2d3a
	13'h169e: q3 = 16'hd6ed; // 0x2d3c
	13'h169f: q3 = 16'h3586; // 0x2d3e
	13'h16a0: q3 = 16'h3a6f; // 0x2d40
	13'h16a1: q3 = 16'hb80a; // 0x2d42
	13'h16a2: q3 = 16'hb59e; // 0x2d44
	13'h16a3: q3 = 16'h192f; // 0x2d46
	13'h16a4: q3 = 16'hc80f; // 0x2d48
	13'h16a5: q3 = 16'h8097; // 0x2d4a
	13'h16a6: q3 = 16'h88e5; // 0x2d4c
	13'h16a7: q3 = 16'hb2c9; // 0x2d4e
	13'h16a8: q3 = 16'h6ed0; // 0x2d50
	13'h16a9: q3 = 16'h0ce3; // 0x2d52
	13'h16aa: q3 = 16'hbf29; // 0x2d54
	13'h16ab: q3 = 16'h40aa; // 0x2d56
	13'h16ac: q3 = 16'hfd65; // 0x2d58
	13'h16ad: q3 = 16'hd720; // 0x2d5a
	13'h16ae: q3 = 16'h3eb2; // 0x2d5c
	13'h16af: q3 = 16'h5d07; // 0x2d5e
	13'h16b0: q3 = 16'hcc0c; // 0x2d60
	13'h16b1: q3 = 16'he594; // 0x2d62
	13'h16b2: q3 = 16'h0d28; // 0x2d64
	13'h16b3: q3 = 16'h8740; // 0x2d66
	13'h16b4: q3 = 16'h219e; // 0x2d68
	13'h16b5: q3 = 16'h1a6e; // 0x2d6a
	13'h16b6: q3 = 16'h001f; // 0x2d6c
	13'h16b7: q3 = 16'h80ba; // 0x2d6e
	13'h16b8: q3 = 16'hf8e8; // 0x2d70
	13'h16b9: q3 = 16'h025a; // 0x2d72
	13'h16ba: q3 = 16'h6e02; // 0x2d74
	13'h16bb: q3 = 16'hd86c; // 0x2d76
	13'h16bc: q3 = 16'h001f; // 0x2d78
	13'h16bd: q3 = 16'h8010; // 0x2d7a
	13'h16be: q3 = 16'h0da5; // 0x2d7c
	13'h16bf: q3 = 16'h86db; // 0x2d7e
	13'h16c0: q3 = 16'hf3b2; // 0x2d80
	13'h16c1: q3 = 16'hf024; // 0x2d82
	13'h16c2: q3 = 16'h940b; // 0x2d84
	13'h16c3: q3 = 16'hb597; // 0x2d86
	13'h16c4: q3 = 16'h6bc0; // 0x2d88
	13'h16c5: q3 = 16'h07e0; // 0x2d8a
	13'h16c6: q3 = 16'h9a1a; // 0x2d8c
	13'h16c7: q3 = 16'h7497; // 0x2d8e
	13'h16c8: q3 = 16'h3036; // 0x2d90
	13'h16c9: q3 = 16'hbe9c; // 0x2d92
	13'h16ca: q3 = 16'h808e; // 0x2d94
	13'h16cb: q3 = 16'h5b21; // 0x2d96
	13'h16cc: q3 = 16'h025b; // 0x2d98
	13'h16cd: q3 = 16'ha3bf; // 0x2d9a
	13'h16ce: q3 = 16'h2940; // 0x2d9c
	13'h16cf: q3 = 16'h07e0; // 0x2d9e
	13'h16d0: q3 = 16'ha6ec; // 0x2da0
	13'h16d1: q3 = 16'hf486; // 0x2da2
	13'h16d2: q3 = 16'hed00; // 0x2da4
	13'h16d3: q3 = 16'hca5c; // 0x2da6
	13'h16d4: q3 = 16'h2c87; // 0x2da8
	13'h16d5: q3 = 16'h9f80; // 0x2daa
	13'h16d6: q3 = 16'hde99; // 0x2dac
	13'h16d7: q3 = 16'h6497; // 0x2dae
	13'h16d8: q3 = 16'h2a2f; // 0x2db0
	13'h16d9: q3 = 16'hb35b; // 0x2db2
	13'h16da: q3 = 16'ha7f8; // 0x2db4
	13'h16db: q3 = 16'hca5c; // 0x2db6
	13'h16dc: q3 = 16'h25d2; // 0x2db8
	13'h16dd: q3 = 16'h98e9; // 0x2dba
	13'h16de: q3 = 16'hbee0; // 0x2dbc
	13'h16df: q3 = 16'h29bb; // 0x2dbe
	13'h16e0: q3 = 16'h3d21; // 0x2dc0
	13'h16e1: q3 = 16'hbb48; // 0x2dc2
	13'h16e2: q3 = 16'h6e96; // 0x2dc4
	13'h16e3: q3 = 16'h1f80; // 0x2dc6
	13'h16e4: q3 = 16'hca5c; // 0x2dc8
	13'h16e5: q3 = 16'h25d2; // 0x2dca
	13'h16e6: q3 = 16'h9d29; // 0x2dcc
	13'h16e7: q3 = 16'hbee0; // 0x2dce
	13'h16e8: q3 = 16'h29bb; // 0x2dd0
	13'h16e9: q3 = 16'h3d21; // 0x2dd2
	13'h16ea: q3 = 16'hbb48; // 0x2dd4
	13'h16eb: q3 = 16'h6e96; // 0x2dd6
	13'h16ec: q3 = 16'h5f80; // 0x2dd8
	13'h16ed: q3 = 16'h961d; // 0x2dda
	13'h16ee: q3 = 16'h00d2; // 0x2ddc
	13'h16ef: q3 = 16'h8940; // 0x2dde
	13'h16f0: q3 = 16'h8efb; // 0x2de0
	13'h16f1: q3 = 16'ha500; // 0x2de2
	13'h16f2: q3 = 16'h1f80; // 0x2de4
	13'h16f3: q3 = 16'hde19; // 0x2de6
	13'h16f4: q3 = 16'ha696; // 0x2de8
	13'h16f5: q3 = 16'hc025; // 0x2dea
	13'h16f6: q3 = 16'hcf39; // 0x2dec
	13'h16f7: q3 = 16'h6e00; // 0x2dee
	13'h16f8: q3 = 16'h1f80; // 0x2df0
	13'h16f9: q3 = 16'h1008; // 0x2df2
	13'h16fa: q3 = 16'hefb6; // 0x2df4
	13'h16fb: q3 = 16'h1ce5; // 0x2df6
	13'h16fc: q3 = 16'h025b; // 0x2df8
	13'h16fd: q3 = 16'h008a; // 0x2dfa
	13'h16fe: q3 = 16'h1cb1; // 0x2dfc
	13'h16ff: q3 = 16'hd69b; // 0x2dfe
	13'h1700: q3 = 16'h2cbc; // 0x2e00
	13'h1701: q3 = 16'h007e; // 0x2e02
	13'h1702: q3 = 16'hb61b; // 0x2e04
	13'h1703: q3 = 16'ha797; // 0x2e06
	13'h1704: q3 = 16'ha02c; // 0x2e08
	13'h1705: q3 = 16'h9408; // 0x2e0a
	13'h1706: q3 = 16'hefca; // 0x2e0c
	13'h1707: q3 = 16'he974; // 0x2e0e
	13'h1708: q3 = 16'h001f; // 0x2e10
	13'h1709: q3 = 16'h80c2; // 0x2e12
	13'h170a: q3 = 16'hc879; // 0x2e14
	13'h170b: q3 = 16'h9720; // 0x2e16
	13'h170c: q3 = 16'h3ecf; // 0x2e18
	13'h170d: q3 = 16'h0a65; // 0x2e1a
	13'h170e: q3 = 16'hb25c; // 0x2e1c
	13'h170f: q3 = 16'h80f8; // 0x2e1e
	13'h1710: q3 = 16'hab59; // 0x2e20
	13'h1711: q3 = 16'he192; // 0x2e22
	13'h1712: q3 = 16'hfc80; // 0x2e24
	13'h1713: q3 = 16'hf8aa; // 0x2e26
	13'h1714: q3 = 16'hfd65; // 0x2e28
	13'h1715: q3 = 16'hd720; // 0x2e2a
	13'h1716: q3 = 16'h3e8a; // 0x2e2c
	13'h1717: q3 = 16'h1ba1; // 0x2e2e
	13'h1718: q3 = 16'hba1c; // 0x2e30
	13'h1719: q3 = 16'hfe8a; // 0x2e32
	13'h171a: q3 = 16'h1ba1; // 0x2e34
	13'h171b: q3 = 16'hba5b; // 0x2e36
	13'h171c: q3 = 16'hbec2; // 0x2e38
	13'h171d: q3 = 16'hc874; // 0x2e3a
	13'h171e: q3 = 16'h86eb; // 0x2e3c
	13'h171f: q3 = 16'hf3f8; // 0x2e3e
	13'h1720: q3 = 16'h8a1b; // 0x2e40
	13'h1721: q3 = 16'ha1ba; // 0x2e42
	13'h1722: q3 = 16'h5cfe; // 0x2e44
	13'h1723: q3 = 16'hc299; // 0x2e46
	13'h1724: q3 = 16'h73f8; // 0x2e48
	13'h1725: q3 = 16'hc21c; // 0x2e4a
	13'h1726: q3 = 16'hf497; // 0x2e4c
	13'h1727: q3 = 16'h496e; // 0x2e4e
	13'h1728: q3 = 16'hf8c2; // 0x2e50
	13'h1729: q3 = 16'h1cf4; // 0x2e52
	13'h172a: q3 = 16'h96c9; // 0x2e54
	13'h172b: q3 = 16'h73f8; // 0x2e56
	13'h172c: q3 = 16'hd21c; // 0x2e58
	13'h172d: q3 = 16'hb497; // 0x2e5a
	13'h172e: q3 = 16'h3f80; // 0x2e5c
	13'h172f: q3 = 16'hc258; // 0x2e5e
	13'h1730: q3 = 16'h73f8; // 0x2e60
	13'h1731: q3 = 16'h9728; // 0x2e62
	13'h1732: q3 = 16'hb396; // 0x2e64
	13'h1733: q3 = 16'hef80; // 0x2e66
	13'h1734: q3 = 16'h9f5a; // 0x2e68
	13'h1735: q3 = 16'h7386; // 0x2e6a
	13'h1736: q3 = 16'hed25; // 0x2e6c
	13'h1737: q3 = 16'hcfe0; // 0x2e6e
	13'h1738: q3 = 16'hc2fa; // 0x2e70
	13'h1739: q3 = 16'h73f8; // 0x2e72
	13'h173a: q3 = 16'hd2fb; // 0x2e74
	13'h173b: q3 = 16'h61d2; // 0x2e76
	13'h173c: q3 = 16'hf973; // 0x2e78
	13'h173d: q3 = 16'hf8d2; // 0x2e7a
	13'h173e: q3 = 16'hfb61; // 0x2e7c
	13'h173f: q3 = 16'hd25b; // 0x2e7e
	13'h1740: q3 = 16'hbed2; // 0x2e80
	13'h1741: q3 = 16'hfb61; // 0x2e82
	13'h1742: q3 = 16'hd25c; // 0x2e84
	13'h1743: q3 = 16'hfed2; // 0x2e86
	13'h1744: q3 = 16'hfb61; // 0x2e88
	13'h1745: q3 = 16'hd25c; // 0x2e8a
	13'h1746: q3 = 16'hfede; // 0x2e8c
	13'h1747: q3 = 16'h1d25; // 0x2e8e
	13'h1748: q3 = 16'hcad9; // 0x2e90
	13'h1749: q3 = 16'h6cbe; // 0x2e92
	13'h174a: q3 = 16'hef80; // 0x2e94
	13'h174b: q3 = 16'hde1c; // 0x2e96
	13'h174c: q3 = 16'hf397; // 0x2e98
	13'h174d: q3 = 16'h2b65; // 0x2e9a
	13'h174e: q3 = 16'hb2fb; // 0x2e9c
	13'h174f: q3 = 16'ha5f8; // 0x2e9e
	13'h1750: q3 = 16'hce1b; // 0x2ea0
	13'h1751: q3 = 16'ha4a6; // 0x2ea2
	13'h1752: q3 = 16'h1f80; // 0x2ea4
	13'h1753: q3 = 16'hc21c; // 0x2ea6
	13'h1754: q3 = 16'hf497; // 0x2ea8
	13'h1755: q3 = 16'h1d65; // 0x2eaa
	13'h1756: q3 = 16'hf8cf; // 0x2eac
	13'h1757: q3 = 16'h4874; // 0x2eae
	13'h1758: q3 = 16'ha73d; // 0x2eb0
	13'h1759: q3 = 16'h298f; // 0x2eb2
	13'h175a: q3 = 16'h3000; // 0x2eb4
	13'h175b: q3 = 16'h030d; // 0x2eb6
	13'h175c: q3 = 16'h73a0; // 0x2eb8
	13'h175d: q3 = 16'h0cf4; // 0x2eba
	13'h175e: q3 = 16'h872d; // 0x2ebc
	13'h175f: q3 = 16'h0044; // 0x2ebe
	13'h1760: q3 = 16'h0d2f; // 0x2ec0
	13'h1761: q3 = 16'h025b; // 0x2ec2
	13'h1762: q3 = 16'ha4f8; // 0x2ec4
	13'h1763: q3 = 16'h03e0; // 0x2ec6
	13'h1764: q3 = 16'hbb5b; // 0x2ec8
	13'h1765: q3 = 16'h6297; // 0x2eca
	13'h1766: q3 = 16'h202f; // 0x2ecc
	13'h1767: q3 = 16'h9809; // 0x2ece
	13'h1768: q3 = 16'he1b6; // 0x2ed0
	13'h1769: q3 = 16'h5cfe; // 0x2ed2
	13'h176a: q3 = 16'h02fb; // 0x2ed4
	13'h176b: q3 = 16'ha537; // 0x2ed6
	13'h176c: q3 = 16'h0b21; // 0x2ed8
	13'h176d: q3 = 16'he65c; // 0x2eda
	13'h176e: q3 = 16'hbe03; // 0x2edc
	13'h176f: q3 = 16'h4def; // 0x2ede
	13'h1770: q3 = 16'h370b; // 0x2ee0
	13'h1771: q3 = 16'h21e6; // 0x2ee2
	13'h1772: q3 = 16'h5cbe; // 0x2ee4
	13'h1773: q3 = 16'h034b; // 0x2ee6
	13'h1774: q3 = 16'hf486; // 0x2ee8
	13'h1775: q3 = 16'hcf80; // 0x2eea
	13'h1776: q3 = 16'h8efa; // 0x2eec
	13'h1777: q3 = 16'h6e02; // 0x2eee
	13'h1778: q3 = 16'h3bf5; // 0x2ef0
	13'h1779: q3 = 16'hbb4f; // 0x2ef2
	13'h177a: q3 = 16'h8003; // 0x2ef4
	13'h177b: q3 = 16'h2a67; // 0x2ef6
	13'h177c: q3 = 16'ha34f; // 0x2ef8
	13'h177d: q3 = 16'h8002; // 0x2efa
	13'h177e: q3 = 16'hc966; // 0x2efc
	13'h177f: q3 = 16'hd3e0; // 0x2efe
	13'h1780: q3 = 16'h8f29; // 0x2f00
	13'h1781: q3 = 16'h64a7; // 0x2f02
	13'h1782: q3 = 16'h4cfe; // 0x2f04
	13'h1783: q3 = 16'h0308; // 0x2f06
	13'h1784: q3 = 16'h6993; // 0x2f08
	13'h1785: q3 = 16'he002; // 0x2f0a
	13'h1786: q3 = 16'h6ca5; // 0x2f0c
	13'h1787: q3 = 16'h97e0; // 0x2f0e
	13'h1788: q3 = 16'h034b; // 0x2f10
	13'h1789: q3 = 16'hf486; // 0x2f12
	13'h178a: q3 = 16'hcf80; // 0x2f14
	13'h178b: q3 = 16'h8afb; // 0x2f16
	13'h178c: q3 = 16'hb5cc; // 0x2f18
	13'h178d: q3 = 16'h0b65; // 0x2f1a
	13'h178e: q3 = 16'hb809; // 0x2f1c
	13'h178f: q3 = 16'h61ca; // 0x2f1e
	13'h1790: q3 = 16'he964; // 0x2f20
	13'h1791: q3 = 16'hf802; // 0x2f22
	13'h1792: q3 = 16'h1d00; // 0x2f24
	13'h1793: q3 = 16'h9a9c; // 0x2f26
	13'h1794: q3 = 16'hb3d0; // 0x2f28
	13'h1795: q3 = 16'h0cf4; // 0x2f2a
	13'h1796: q3 = 16'h8679; // 0x2f2c
	13'h1797: q3 = 16'h7e02; // 0x2f2e
	13'h1798: q3 = 16'h1d00; // 0x2f30
	13'h1799: q3 = 16'ha299; // 0x2f32
	13'h179a: q3 = 16'he897; // 0x2f34
	13'h179b: q3 = 16'h2033; // 0x2f36
	13'h179c: q3 = 16'hd219; // 0x2f38
	13'h179d: q3 = 16'he5cf; // 0x2f3a
	13'h179e: q3 = 16'he003; // 0x2f3c
	13'h179f: q3 = 16'h7a74; // 0x2f3e
	13'h17a0: q3 = 16'ha00b; // 0x2f40
	13'h17a1: q3 = 16'h25da; // 0x2f42
	13'h17a2: q3 = 16'h5b00; // 0x2f44
	13'h17a3: q3 = 16'hce5b; // 0x2f46
	13'h17a4: q3 = 16'h258f; // 0x2f48
	13'h17a5: q3 = 16'h4f80; // 0x2f4a
	13'h17a6: q3 = 16'h034b; // 0x2f4c
	13'h17a7: q3 = 16'hf486; // 0x2f4e
	13'h17a8: q3 = 16'hcf80; // 0x2f50
	13'h17a9: q3 = 16'h0278; // 0x2f52
	13'h17aa: q3 = 16'h6d97; // 0x2f54
	13'h17ab: q3 = 16'h3037; // 0x2f56
	13'h17ac: q3 = 16'ha74a; // 0x2f58
	13'h17ad: q3 = 16'h008a; // 0x2f5a
	13'h17ae: q3 = 16'hfbb5; // 0x2f5c
	13'h17af: q3 = 16'hcc0b; // 0x2f5e
	13'h17b0: q3 = 16'h65bb; // 0x2f60
	13'h17b1: q3 = 16'he087; // 0x2f62
	13'h17b2: q3 = 16'h6972; // 0x2f64
	13'h17b3: q3 = 16'h8679; // 0x2f66
	13'h17b4: q3 = 16'h40d2; // 0x2f68
	13'h17b5: q3 = 16'h9b65; // 0x2f6a
	13'h17b6: q3 = 16'hf802; // 0x2f6c
	13'h17b7: q3 = 16'h2974; // 0x2f6e
	13'h17b8: q3 = 16'hde59; // 0x2f70
	13'h17b9: q3 = 16'h6e02; // 0x2f72
	13'h17ba: q3 = 16'h3ca5; // 0x2f74
	13'h17bb: q3 = 16'h929d; // 0x2f76
	13'h17bc: q3 = 16'h33f8; // 0x2f78
	13'h17bd: q3 = 16'h0309; // 0x2f7a
	13'h17be: q3 = 16'h7202; // 0x2f7c
	13'h17bf: q3 = 16'h786d; // 0x2f7e
	13'h17c0: q3 = 16'h97e0; // 0x2f80
	13'h17c1: q3 = 16'hb2fb; // 0x2f82
	13'h17c2: q3 = 16'ha702; // 0x2f84
	13'h17c3: q3 = 16'h786d; // 0x2f86
	13'h17c4: q3 = 16'h97e0; // 0x2f88
	13'h17c5: q3 = 16'hd2fd; // 0x2f8a
	13'h17c6: q3 = 16'h21b0; // 0x2f8c
	13'h17c7: q3 = 16'h0d29; // 0x2f8e
	13'h17c8: q3 = 16'hb650; // 0x2f90
	13'h17c9: q3 = 16'h2fbb; // 0x2f92
	13'h17ca: q3 = 16'he0a6; // 0x2f94
	13'h17cb: q3 = 16'he030; // 0x2f96
	13'h17cc: q3 = 16'hb21e; // 0x2f98
	13'h17cd: q3 = 16'h40b6; // 0x2f9a
	13'h17ce: q3 = 16'hf925; // 0x2f9c
	13'h17cf: q3 = 16'hf803; // 0x2f9e
	13'h17d0: q3 = 16'he0d2; // 0x2fa0
	13'h17d1: q3 = 16'hfd21; // 0x2fa2
	13'h17d2: q3 = 16'hb00d; // 0x2fa4
	13'h17d3: q3 = 16'h29b6; // 0x2fa6
	13'h17d4: q3 = 16'h5f80; // 0x2fa8
	13'h17d5: q3 = 16'hd2fd; // 0x2faa
	13'h17d6: q3 = 16'h21b0; // 0x2fac
	13'h17d7: q3 = 16'h08f2; // 0x2fae
	13'h17d8: q3 = 16'h964a; // 0x2fb0
	13'h17d9: q3 = 16'h74cc; // 0x2fb2
	13'h17da: q3 = 16'h0000; // 0x2fb4
	13'h17db: q3 = 16'h0000; // 0x2fb6
	13'h17dc: q3 = 16'h0000; // 0x2fb8
	13'h17dd: q3 = 16'h0000; // 0x2fba
	13'h17de: q3 = 16'h000f; // 0x2fbc
	13'h17df: q3 = 16'h80d2; // 0x2fbe
	13'h17e0: q3 = 16'h5cf4; // 0x2fc0
	13'h17e1: q3 = 16'hcfe0; // 0x2fc2
	13'h17e2: q3 = 16'hcf48; // 0x2fc4
	13'h17e3: q3 = 16'h74a7; // 0x2fc6
	13'h17e4: q3 = 16'h3d29; // 0x2fc8
	13'h17e5: q3 = 16'h8f3f; // 0x2fca
	13'h17e6: q3 = 16'h80bf; // 0x2fcc
	13'h17e7: q3 = 16'h0d29; // 0x2fce
	13'h17e8: q3 = 16'hbeec; // 0x2fd0
	13'h17e9: q3 = 16'hfece; // 0x2fd2
	13'h17ea: q3 = 16'h5b26; // 0x2fd4
	13'h17eb: q3 = 16'h3749; // 0x2fd6
	13'h17ec: q3 = 16'h73d3; // 0x2fd8
	13'h17ed: q3 = 16'he0b6; // 0x2fda
	13'h17ee: q3 = 16'hfda5; // 0x2fdc
	13'h17ef: q3 = 16'h02ab; // 0x2fde
	13'h17f0: q3 = 16'hf9cf; // 0x2fe0
	13'h17f1: q3 = 16'h4a63; // 0x2fe2
	13'h17f2: q3 = 16'hac0d; // 0x2fe4
	13'h17f3: q3 = 16'h2f02; // 0x2fe6
	13'h17f4: q3 = 16'h3a21; // 0x2fe8
	13'h17f5: q3 = 16'hba79; // 0x2fea
	13'h17f6: q3 = 16'h7ec3; // 0x2fec
	13'h17f7: q3 = 16'h5ce8; // 0x2fee
	13'h17f8: q3 = 16'h034a; // 0x2ff0
	13'h17f9: q3 = 16'h32bf; // 0x2ff2
	13'h17fa: q3 = 16'h7034; // 0x2ff4
	13'h17fb: q3 = 16'hbc0c; // 0x2ff6
	13'h17fc: q3 = 16'he5b2; // 0x2ff8
	13'h17fd: q3 = 16'h58f4; // 0x2ffa
	13'h17fe: q3 = 16'hf8d3; // 0x2ffc
	13'h17ff: q3 = 16'h5cae; // 0x2ffe
	13'h1800: q3 = 16'h0339; // 0x3000
	13'h1801: q3 = 16'h6c98; // 0x3002
	13'h1802: q3 = 16'hdd25; // 0x3004
	13'h1803: q3 = 16'hcf40; // 0x3006
	13'h1804: q3 = 16'h33de; // 0x3008
	13'h1805: q3 = 16'h9d23; // 0x300a
	13'h1806: q3 = 16'ha00b; // 0x300c
	13'h1807: q3 = 16'he698; // 0x300e
	13'h1808: q3 = 16'h0d2f; // 0x3010
	13'h1809: q3 = 16'h025b; // 0x3012
	13'h180a: q3 = 16'ha4f8; // 0x3014
	13'h180b: q3 = 16'haafe; // 0x3016
	13'h180c: q3 = 16'h73d2; // 0x3018
	13'h180d: q3 = 16'h98eb; // 0x301a
	13'h180e: q3 = 16'h0238; // 0x301c
	13'h180f: q3 = 16'h6ca6; // 0x301e
	13'h1810: q3 = 16'h2ca1; // 0x3020
	13'h1811: q3 = 16'hd29b; // 0x3022
	13'h1812: q3 = 16'heef8; // 0x3024
	13'h1813: q3 = 16'hcf7a; // 0x3026
	13'h1814: q3 = 16'h748e; // 0x3028
	13'h1815: q3 = 16'h8034; // 0x302a
	13'h1816: q3 = 16'h973d; // 0x302c
	13'h1817: q3 = 16'h3e8e; // 0x302e
	13'h1818: q3 = 16'hfb2f; // 0x3030
	13'h1819: q3 = 16'hc80c; // 0x3032
	13'h181a: q3 = 16'h21d3; // 0x3034
	13'h181b: q3 = 16'h4972; // 0x3036
	13'h181c: q3 = 16'hbbe0; // 0x3038
	13'h181d: q3 = 16'h8efb; // 0x303a
	13'h181e: q3 = 16'hb697; // 0x303c
	13'h181f: q3 = 16'h29e5; // 0x303e
	13'h1820: q3 = 16'hba39; // 0x3040
	13'h1821: q3 = 16'h40c2; // 0x3042
	13'h1822: q3 = 16'h1d34; // 0x3044
	13'h1823: q3 = 16'h972b; // 0x3046
	13'h1824: q3 = 16'hbece; // 0x3048
	13'h1825: q3 = 16'hfd6e; // 0x304a
	13'h1826: q3 = 16'h900d; // 0x304c
	13'h1827: q3 = 16'h25cf; // 0x304e
	13'h1828: q3 = 16'h4f80; // 0x3050
	13'h1829: q3 = 16'hd25c; // 0x3052
	13'h182a: q3 = 16'hf4cf; // 0x3054
	13'h182b: q3 = 16'he0c3; // 0x3056
	13'h182c: q3 = 16'h5ce8; // 0x3058
	13'h182d: q3 = 16'h033d; // 0x305a
	13'h182e: q3 = 16'h21cb; // 0x305c
	13'h182f: q3 = 16'h4011; // 0x305e
	13'h1830: q3 = 16'h034b; // 0x3060
	13'h1831: q3 = 16'hc096; // 0x3062
	13'h1832: q3 = 16'he900; // 0x3064
	13'h1833: q3 = 16'hd25c; // 0x3066
	13'h1834: q3 = 16'hf4cf; // 0x3068
	13'h1835: q3 = 16'he0aa; // 0x306a
	13'h1836: q3 = 16'hfe73; // 0x306c
	13'h1837: q3 = 16'hd298; // 0x306e
	13'h1838: q3 = 16'heb02; // 0x3070
	13'h1839: q3 = 16'h386c; // 0x3072
	13'h183a: q3 = 16'ha62c; // 0x3074
	13'h183b: q3 = 16'ha1d2; // 0x3076
	13'h183c: q3 = 16'h9bee; // 0x3078
	13'h183d: q3 = 16'hf8a2; // 0x307a
	13'h183e: q3 = 16'hfb24; // 0x307c
	13'h183f: q3 = 16'h02ab; // 0x307e
	13'h1840: q3 = 16'hf9cf; // 0x3080
	13'h1841: q3 = 16'h4a63; // 0x3082
	13'h1842: q3 = 16'hac0a; // 0x3084
	13'h1843: q3 = 16'h6e02; // 0x3086
	13'h1844: q3 = 16'h5863; // 0x3088
	13'h1845: q3 = 16'ha009; // 0x308a
	13'h1846: q3 = 16'h29ca; // 0x308c
	13'h1847: q3 = 16'h58f4; // 0x308e
	13'h1848: q3 = 16'ha6fb; // 0x3090
	13'h1849: q3 = 16'hbe9a; // 0x3092
	13'h184a: q3 = 16'hfc80; // 0x3094
	13'h184b: q3 = 16'h9a9d; // 0x3096
	13'h184c: q3 = 16'ha503; // 0x3098
	13'h184d: q3 = 16'h3963; // 0x309a
	13'h184e: q3 = 16'hbee9; // 0x309c
	13'h184f: q3 = 16'h33f8; // 0x309e
	13'h1850: q3 = 16'hc35c; // 0x30a0
	13'h1851: q3 = 16'he803; // 0x30a2
	13'h1852: q3 = 16'h3d21; // 0x30a4
	13'h1853: q3 = 16'hcb40; // 0x30a6
	13'h1854: q3 = 16'h1203; // 0x30a8
	13'h1855: q3 = 16'h4bc0; // 0x30aa
	13'h1856: q3 = 16'h8e1b; // 0x30ac
	13'h1857: q3 = 16'h298b; // 0x30ae
	13'h1858: q3 = 16'h2874; // 0x30b0
	13'h1859: q3 = 16'h97e0; // 0x30b2
	13'h185a: q3 = 16'hc2c8; // 0x30b4
	13'h185b: q3 = 16'h7997; // 0x30b6
	13'h185c: q3 = 16'h2000; // 0x30b8
	13'h185d: q3 = 16'h02ab; // 0x30ba
	13'h185e: q3 = 16'hf9cf; // 0x30bc
	13'h185f: q3 = 16'h4a63; // 0x30be
	13'h1860: q3 = 16'hafe0; // 0x30c0
	13'h1861: q3 = 16'hc35c; // 0x30c2
	13'h1862: q3 = 16'he803; // 0x30c4
	13'h1863: q3 = 16'h3d21; // 0x30c6
	13'h1864: q3 = 16'hcb40; // 0x30c8
	13'h1865: q3 = 16'h1103; // 0x30ca
	13'h1866: q3 = 16'h4bc0; // 0x30cc
	13'h1867: q3 = 16'h96e9; // 0x30ce
	13'h1868: q3 = 16'h3ece; // 0x30d0
	13'h1869: q3 = 16'hfd6e; // 0x30d2
	13'h186a: q3 = 16'h900d; // 0x30d4
	13'h186b: q3 = 16'h25cf; // 0x30d6
	13'h186c: q3 = 16'h4f80; // 0x30d8
	13'h186d: q3 = 16'h8e88; // 0x30da
	13'h186e: q3 = 16'h6eba; // 0x30dc
	13'h186f: q3 = 16'h5b00; // 0x30de
	13'h1870: q3 = 16'h000f; // 0x30e0
	13'h1871: q3 = 16'h80c3; // 0x30e2
	13'h1872: q3 = 16'h5ce8; // 0x30e4
	13'h1873: q3 = 16'h033d; // 0x30e6
	13'h1874: q3 = 16'h21cb; // 0x30e8
	13'h1875: q3 = 16'h4011; // 0x30ea
	13'h1876: q3 = 16'h034b; // 0x30ec
	13'h1877: q3 = 16'hc096; // 0x30ee
	13'h1878: q3 = 16'he93e; // 0x30f0
	13'h1879: q3 = 16'hcf7a; // 0x30f2
	13'h187a: q3 = 16'h748e; // 0x30f4
	13'h187b: q3 = 16'h8034; // 0x30f6
	13'h187c: q3 = 16'h973d; // 0x30f8
	13'h187d: q3 = 16'h3ec3; // 0x30fa
	13'h187e: q3 = 16'h5ce8; // 0x30fc
	13'h187f: q3 = 16'h033d; // 0x30fe
	13'h1880: q3 = 16'h21cb; // 0x3100
	13'h1881: q3 = 16'h4011; // 0x3102
	13'h1882: q3 = 16'h021b; // 0x3104
	13'h1883: q3 = 16'ha403; // 0x3106
	13'h1884: q3 = 16'h3d21; // 0x3108
	13'h1885: q3 = 16'hcb40; // 0x310a
	13'h1886: q3 = 16'h1203; // 0x310c
	13'h1887: q3 = 16'h4bc0; // 0x310e
	13'h1888: q3 = 16'h96e9; // 0x3110
	13'h1889: q3 = 16'h3ecf; // 0x3112
	13'h188a: q3 = 16'h4872; // 0x3114
	13'h188b: q3 = 16'hd004; // 0x3116
	13'h188c: q3 = 16'h7ecf; // 0x3118
	13'h188d: q3 = 16'h4872; // 0x311a
	13'h188e: q3 = 16'hd004; // 0x311c
	13'h188f: q3 = 16'hbed2; // 0x311e
	13'h1890: q3 = 16'h8caf; // 0x3120
	13'h1891: q3 = 16'hdc04; // 0x3122
	13'h1892: q3 = 16'h7eaa; // 0x3124
	13'h1893: q3 = 16'hfe73; // 0x3126
	13'h1894: q3 = 16'hd298; // 0x3128
	13'h1895: q3 = 16'heb01; // 0x312a
	13'h1896: q3 = 16'h1f80; // 0x312c
	13'h1897: q3 = 16'h000e; // 0x312e
	13'h1898: q3 = 16'h3e00; // 0x3130
	13'h1899: q3 = 16'h0e7e; // 0x3132
	13'h189a: q3 = 16'hb259; // 0x3134
	13'h189b: q3 = 16'hb402; // 0x3136
	13'h189c: q3 = 16'h3be9; // 0x3138
	13'h189d: q3 = 16'hbbe0; // 0x313a
	13'h189e: q3 = 16'hca99; // 0x313c
	13'h189f: q3 = 16'he8d0; // 0x313e
	13'h18a0: q3 = 16'h08ef; // 0x3140
	13'h18a1: q3 = 16'ha6ef; // 0x3142
	13'h18a2: q3 = 16'h8087; // 0x3144
	13'h18a3: q3 = 16'h5e00; // 0x3146
	13'h18a4: q3 = 16'h8efa; // 0x3148
	13'h18a5: q3 = 16'h6ef8; // 0x314a
	13'h18a6: q3 = 16'h929c; // 0x314c
	13'h18a7: q3 = 16'h00cf; // 0x314e
	13'h18a8: q3 = 16'h7a74; // 0x3150
	13'h18a9: q3 = 16'h8e89; // 0x3152
	13'h18aa: q3 = 16'h7300; // 0x3154
	13'h18ab: q3 = 16'h0011; // 0x3156
	13'h18ac: q3 = 16'h0120; // 0x3158
	13'h18ad: q3 = 16'h1301; // 0x315a
	13'h18ae: q3 = 16'h4015; // 0x315c
	13'h18af: q3 = 16'h0160; // 0x315e
	13'h18b0: q3 = 16'h1701; // 0x3160
	13'h18b1: q3 = 16'h8f80; // 0x3162
	13'h18b2: q3 = 16'hd28c; // 0x3164
	13'h18b3: q3 = 16'hafdc; // 0x3166
	13'h18b4: q3 = 16'h04be; // 0x3168
	13'h18b5: q3 = 16'haafe; // 0x316a
	13'h18b6: q3 = 16'h73d2; // 0x316c
	13'h18b7: q3 = 16'h98eb; // 0x316e
	13'h18b8: q3 = 16'h012f; // 0x3170
	13'h18b9: q3 = 16'h8000; // 0x3172
	13'h18ba: q3 = 16'h0e3e; // 0x3174
	13'h18bb: q3 = 16'h000e; // 0x3176
	13'h18bc: q3 = 16'h7ebf; // 0x3178
	13'h18bd: q3 = 16'h0d29; // 0x317a
	13'h18be: q3 = 16'hbeec; // 0x317c
	13'h18bf: q3 = 16'hfeb6; // 0x317e
	13'h18c0: q3 = 16'hfda5; // 0x3180
	13'h18c1: q3 = 16'h02ab; // 0x3182
	13'h18c2: q3 = 16'hf9cf; // 0x3184
	13'h18c3: q3 = 16'h4a63; // 0x3186
	13'h18c4: q3 = 16'hac0d; // 0x3188
	13'h18c5: q3 = 16'h2f02; // 0x318a
	13'h18c6: q3 = 16'h3a21; // 0x318c
	13'h18c7: q3 = 16'hba79; // 0x318e
	13'h18c8: q3 = 16'h40ca; // 0x3190
	13'h18c9: q3 = 16'hfdfe; // 0x3192
	13'h18ca: q3 = 16'hc35c; // 0x3194
	13'h18cb: q3 = 16'he803; // 0x3196
	13'h18cc: q3 = 16'h4a32; // 0x3198
	13'h18cd: q3 = 16'hbf70; // 0x319a
	13'h18ce: q3 = 16'h34bc; // 0x319c
	13'h18cf: q3 = 16'h08e8; // 0x319e
	13'h18d0: q3 = 16'h86e9; // 0x31a0
	13'h18d1: q3 = 16'he503; // 0x31a2
	13'h18d2: q3 = 16'h3974; // 0x31a4
	13'h18d3: q3 = 16'hd29b; // 0x31a6
	13'h18d4: q3 = 16'ha7cf; // 0x31a8
	13'h18d5: q3 = 16'he0c3; // 0x31aa
	13'h18d6: q3 = 16'h5ce8; // 0x31ac
	13'h18d7: q3 = 16'h033d; // 0x31ae
	13'h18d8: q3 = 16'h21cb; // 0x31b0
	13'h18d9: q3 = 16'h4011; // 0x31b2
	13'h18da: q3 = 16'h034b; // 0x31b4
	13'h18db: q3 = 16'hc096; // 0x31b6
	13'h18dc: q3 = 16'he93e; // 0x31b8
	13'h18dd: q3 = 16'hce5d; // 0x31ba
	13'h18de: q3 = 16'h34a6; // 0x31bc
	13'h18df: q3 = 16'he9f3; // 0x31be
	13'h18e0: q3 = 16'hf8ca; // 0x31c0
	13'h18e1: q3 = 16'h5cf4; // 0x31c2
	13'h18e2: q3 = 16'hbf29; // 0x31c4
	13'h18e3: q3 = 16'h40ce; // 0x31c6
	13'h18e4: q3 = 16'h5d34; // 0x31c8
	13'h18e5: q3 = 16'ha6e9; // 0x31ca
	13'h18e6: q3 = 16'hf3f8; // 0x31cc
	13'h18e7: q3 = 16'h8ec9; // 0x31ce
	13'h18e8: q3 = 16'h61c8; // 0x31d0
	13'h18e9: q3 = 16'h0da1; // 0x31d2
	13'h18ea: q3 = 16'hb359; // 0x31d4
	13'h18eb: q3 = 16'h73f8; // 0x31d6
	13'h18ec: q3 = 16'hb29d; // 0x31d8
	13'h18ed: q3 = 16'ha5cc; // 0x31da
	13'h18ee: q3 = 16'h0c25; // 0x31dc
	13'h18ef: q3 = 16'hc809; // 0x31de
	13'h18f0: q3 = 16'he1b6; // 0x31e0
	13'h18f1: q3 = 16'h5f80; // 0x31e2
	13'h18f2: q3 = 16'h9299; // 0x31e4
	13'h18f3: q3 = 16'ha6a6; // 0x31e6
	13'h18f4: q3 = 16'h3d6c; // 0x31e8
	13'h18f5: q3 = 16'hd39f; // 0x31ea
	13'h18f6: q3 = 16'h809a; // 0x31ec
	13'h18f7: q3 = 16'h9cb3; // 0x31ee
	13'h18f8: q3 = 16'hd008; // 0x31f0
	13'h18f9: q3 = 16'hafbb; // 0x31f2
	13'h18fa: q3 = 16'h5cc0; // 0x31f4
	13'h18fb: q3 = 16'hcf48; // 0x31f6
	13'h18fc: q3 = 16'h6797; // 0x31f8
	13'h18fd: q3 = 16'he0a2; // 0x31fa
	13'h18fe: q3 = 16'h99e8; // 0x31fc
	13'h18ff: q3 = 16'h9720; // 0x31fe
	13'h1900: q3 = 16'h22be; // 0x3200
	13'h1901: q3 = 16'hed73; // 0x3202
	13'h1902: q3 = 16'h033d; // 0x3204
	13'h1903: q3 = 16'h219e; // 0x3206
	13'h1904: q3 = 16'h5f80; // 0x3208
	13'h1905: q3 = 16'hb25d; // 0x320a
	13'h1906: q3 = 16'ha5b0; // 0x320c
	13'h1907: q3 = 16'h0ce5; // 0x320e
	13'h1908: q3 = 16'hb258; // 0x3210
	13'h1909: q3 = 16'hf402; // 0x3212
	13'h190a: q3 = 16'h2bee; // 0x3214
	13'h190b: q3 = 16'hd73f; // 0x3216
	13'h190c: q3 = 16'h80b2; // 0x3218
	13'h190d: q3 = 16'h5da5; // 0x321a
	13'h190e: q3 = 16'hb00c; // 0x321c
	13'h190f: q3 = 16'he5b2; // 0x321e
	13'h1910: q3 = 16'h58f4; // 0x3220
	13'h1911: q3 = 16'h02db; // 0x3222
	13'h1912: q3 = 16'he497; // 0x3224
	13'h1913: q3 = 16'he087; // 0x3226
	13'h1914: q3 = 16'h4d32; // 0x3228
	13'h1915: q3 = 16'h863d; // 0x322a
	13'h1916: q3 = 16'h00ce; // 0x322c
	13'h1917: q3 = 16'hfd6e; // 0x322e
	13'h1918: q3 = 16'h933f; // 0x3230
	13'h1919: q3 = 16'h80b2; // 0x3232
	13'h191a: q3 = 16'h1ba7; // 0x3234
	13'h191b: q3 = 16'hd619; // 0x3236
	13'h191c: q3 = 16'he5f8; // 0x3238
	13'h191d: q3 = 16'h8ef8; // 0x323a
	13'h191e: q3 = 16'hebd2; // 0x323c
	13'h191f: q3 = 16'h1a6c; // 0x323e
	13'h1920: q3 = 16'h02db; // 0x3240
	13'h1921: q3 = 16'he497; // 0x3242
	13'h1922: q3 = 16'he08e; // 0x3244
	13'h1923: q3 = 16'hfa6e; // 0x3246
	13'h1924: q3 = 16'h023b; // 0x3248
	13'h1925: q3 = 16'hf5bb; // 0x324a
	13'h1926: q3 = 16'h4972; // 0x324c
	13'h1927: q3 = 16'hcfe0; // 0x324e
	13'h1928: q3 = 16'h8f5c; // 0x3250
	13'h1929: q3 = 16'hb296; // 0x3252
	13'h192a: q3 = 16'hed3e; // 0x3254
	13'h192b: q3 = 16'h9a18; // 0x3256
	13'h192c: q3 = 16'hf4bf; // 0x3258
	13'h192d: q3 = 16'h2e7e; // 0x325a
	13'h192e: q3 = 16'ha299; // 0x325c
	13'h192f: q3 = 16'he803; // 0x325e
	13'h1930: q3 = 16'h38ef; // 0x3260
	13'h1931: q3 = 16'hca5c; // 0x3262
	13'h1932: q3 = 16'hfecf; // 0x3264
	13'h1933: q3 = 16'h4874; // 0x3266
	13'h1934: q3 = 16'ha73d; // 0x3268
	13'h1935: q3 = 16'h298f; // 0x326a
	13'h1936: q3 = 16'h3f80; // 0x326c
	13'h1937: q3 = 16'h47e0; // 0x326e
	13'h1938: q3 = 16'h4be0; // 0x3270
	13'h1939: q3 = 16'h4fe0; // 0x3272
	13'h193a: q3 = 16'h53e0; // 0x3274
	13'h193b: q3 = 16'h57e0; // 0x3276
	13'h193c: q3 = 16'hbe69; // 0x3278
	13'h193d: q3 = 16'hbebe; // 0x327a
	13'h193e: q3 = 16'hef80; // 0x327c
	13'h193f: q3 = 16'hbafc; // 0x327e
	13'h1940: q3 = 16'had86; // 0x3280
	13'h1941: q3 = 16'hcf80; // 0x3282
	13'h1942: q3 = 16'h8efb; // 0x3284
	13'h1943: q3 = 16'hb3d2; // 0x3286
	13'h1944: q3 = 16'h1bb4; // 0x3288
	13'h1945: q3 = 16'hf892; // 0x328a
	13'h1946: q3 = 16'h5b6f; // 0x328c
	13'h1947: q3 = 16'hf8be; // 0x328e
	13'h1948: q3 = 16'h69be; // 0x3290
	13'h1949: q3 = 16'h96e9; // 0x3292
	13'h194a: q3 = 16'heca7; // 0x3294
	13'h194b: q3 = 16'h3a3e; // 0x3296
	13'h194c: q3 = 16'h9e5c; // 0x3298
	13'h194d: q3 = 16'had86; // 0x329a
	13'h194e: q3 = 16'hef80; // 0x329c
	13'h194f: q3 = 16'hcf08; // 0x329e
	13'h1950: q3 = 16'h6ea7; // 0x32a0
	13'h1951: q3 = 16'h3a3e; // 0x32a2
	13'h1952: q3 = 16'h9b29; // 0x32a4
	13'h1953: q3 = 16'h6e8e; // 0x32a6
	13'h1954: q3 = 16'h8f80; // 0x32a8
	13'h1955: q3 = 16'hbee9; // 0x32aa
	13'h1956: q3 = 16'h7ed3; // 0x32ac
	13'h1957: q3 = 16'h7bfe; // 0x32ae
	13'h1958: q3 = 16'h03e0; // 0x32b0
	13'h1959: q3 = 16'hc35c; // 0x32b2
	13'h195a: q3 = 16'he803; // 0x32b4
	13'h195b: q3 = 16'h4a32; // 0x32b6
	13'h195c: q3 = 16'hbf7f; // 0x32b8
	13'h195d: q3 = 16'h80ca; // 0x32ba
	13'h195e: q3 = 16'h5cf4; // 0x32bc
	13'h195f: q3 = 16'hbf29; // 0x32be
	13'h1960: q3 = 16'h64f8; // 0x32c0
	13'h1961: q3 = 16'h03e0; // 0x32c2
	13'h1962: q3 = 16'hc35c; // 0x32c4
	13'h1963: q3 = 16'he803; // 0x32c6
	13'h1964: q3 = 16'h4a32; // 0x32c8
	13'h1965: q3 = 16'hbf7f; // 0x32ca
	13'h1966: q3 = 16'h808e; // 0x32cc
	13'h1967: q3 = 16'hc961; // 0x32ce
	13'h1968: q3 = 16'hca59; // 0x32d0
	13'h1969: q3 = 16'h3ecf; // 0x32d2
	13'h196a: q3 = 16'h4874; // 0x32d4
	13'h196b: q3 = 16'ha73d; // 0x32d6
	13'h196c: q3 = 16'h298f; // 0x32d8
	13'h196d: q3 = 16'h3f80; // 0x32da
	13'h196e: q3 = 16'hd29b; // 0x32dc
	13'h196f: q3 = 16'h6500; // 0x32de
	13'h1970: q3 = 16'h6023; // 0x32e0
	13'h1971: q3 = 16'hca59; // 0x32e2
	13'h1972: q3 = 16'h29d3; // 0x32e4
	13'h1973: q3 = 16'h3f80; // 0x32e6
	13'h1974: q3 = 16'ha299; // 0x32e8
	13'h1975: q3 = 16'he803; // 0x32ea
	13'h1976: q3 = 16'h38ef; // 0x32ec
	13'h1977: q3 = 16'hca5c; // 0x32ee
	13'h1978: q3 = 16'hfebf; // 0x32f0
	13'h1979: q3 = 16'h0d29; // 0x32f2
	13'h197a: q3 = 16'hbeec; // 0x32f4
	13'h197b: q3 = 16'hfeaa; // 0x32f6
	13'h197c: q3 = 16'hfe73; // 0x32f8
	13'h197d: q3 = 16'hd298; // 0x32fa
	13'h197e: q3 = 16'heb03; // 0x32fc
	13'h197f: q3 = 16'h686c; // 0x32fe
	13'h1980: q3 = 16'hd65c; // 0x3300
	13'h1981: q3 = 16'hfebb; // 0x3302
	13'h1982: q3 = 16'h6ca1; // 0x3304
	13'h1983: q3 = 16'hb409; // 0x3306
	13'h1984: q3 = 16'ha1a6; // 0x3308
	13'h1985: q3 = 16'hc964; // 0x330a
	13'h1986: q3 = 16'h6be0; // 0x330c
	13'h1987: q3 = 16'hbb6c; // 0x330e
	13'h1988: q3 = 16'ha1b4; // 0x3310
	13'h1989: q3 = 16'h0beb; // 0x3312
	13'h198a: q3 = 16'hf800; // 0x3314
	13'h198b: q3 = 16'h8000; // 0x3316
	13'h198c: q3 = 16'h0000; // 0x3318
	13'h198d: q3 = 16'h0180; // 0x331a
	13'h198e: q3 = 16'h0180; // 0x331c
	13'h198f: q3 = 16'h0005; // 0x331e
	13'h1990: q3 = 16'h0000; // 0x3320
	13'h1991: q3 = 16'h0000; // 0x3322
	13'h1992: q3 = 16'h000f; // 0x3324
	13'h1993: q3 = 16'hffc0; // 0x3326
	13'h1994: q3 = 16'hffc0; // 0x3328
	13'h1995: q3 = 16'h000e; // 0x332a
	13'h1996: q3 = 16'h0000; // 0x332c
	13'h1997: q3 = 16'h0000; // 0x332e
	13'h1998: q3 = 16'h7fff; // 0x3330
	13'h1999: q3 = 16'h0000; // 0x3332
	13'h199a: q3 = 16'h8136; // 0x3334
	13'h199b: q3 = 16'h0000; // 0x3336
	13'h199c: q3 = 16'hf31a; // 0x3338
	13'h199d: q3 = 16'h0000; // 0x333a
	13'h199e: q3 = 16'h0001; // 0x333c
	13'h199f: q3 = 16'hffd4; // 0x333e
	13'h19a0: q3 = 16'hffec; // 0x3340
	13'h19a1: q3 = 16'h0032; // 0x3342
	13'h19a2: q3 = 16'h0000; // 0x3344
	13'h19a3: q3 = 16'h0000; // 0x3346
	13'h19a4: q3 = 16'h7fff; // 0x3348
	13'h19a5: q3 = 16'h0000; // 0x334a
	13'h19a6: q3 = 16'h8136; // 0x334c
	13'h19a7: q3 = 16'h0000; // 0x334e
	13'h19a8: q3 = 16'hf33e; // 0x3350
	13'h19a9: q3 = 16'h0400; // 0x3352
	13'h19aa: q3 = 16'h0000; // 0x3354
	13'h19ab: q3 = 16'h001f; // 0x3356
	13'h19ac: q3 = 16'h3f7f; // 0x3358
	13'h19ad: q3 = 16'h7f7f; // 0x335a
	13'h19ae: q3 = 16'h7e3f; // 0x335c
	13'h19af: q3 = 16'h1f1f; // 0x335e
	13'h19b0: q3 = 16'h1e1c; // 0x3360
	13'h19b1: q3 = 16'h001f; // 0x3362
	13'h19b2: q3 = 16'h3f7c; // 0x3364
	13'h19b3: q3 = 16'h7f7f; // 0x3366
	13'h19b4: q3 = 16'h7f3f; // 0x3368
	13'h19b5: q3 = 16'h3f1f; // 0x336a
	13'h19b6: q3 = 16'h1f1f; // 0x336c
	13'h19b7: q3 = 16'h3e3f; // 0x336e
	13'h19b8: q3 = 16'h3f3e; // 0x3370
	13'h19b9: q3 = 16'h3830; // 0x3372
	13'h19ba: q3 = 16'h3000; // 0x3374
	13'h19bb: q3 = 16'h0d00; // 0x3376
	13'h19bc: q3 = 16'h0000; // 0x3378
	13'h19bd: q3 = 16'hf386; // 0x337a
	13'h19be: q3 = 16'h0d00; // 0x337c
	13'h19bf: q3 = 16'h0000; // 0x337e
	13'h19c0: q3 = 16'hf414; // 0x3380
	13'h19c1: q3 = 16'h0801; // 0x3382
	13'h19c2: q3 = 16'h0100; // 0x3384
	13'h19c3: q3 = 16'h0001; // 0x3386
	13'h19c4: q3 = 16'h0200; // 0x3388
	13'h19c5: q3 = 16'h0049; // 0x338a
	13'h19c6: q3 = 16'hf49f; // 0x338c
	13'h19c7: q3 = 16'h0301; // 0x338e
	13'h19c8: q3 = 16'h0000; // 0x3390
	13'h19c9: q3 = 16'hc36e; // 0x3392
	13'h19ca: q3 = 16'h0501; // 0x3394
	13'h19cb: q3 = 16'h0000; // 0x3396
	13'h19cc: q3 = 16'hc386; // 0x3398
	13'h19cd: q3 = 16'h8701; // 0x339a
	13'h19ce: q3 = 16'h0333; // 0x339c
	13'h19cf: q3 = 16'h0666; // 0x339e
	13'h19d0: q3 = 16'h8a01; // 0x33a0
	13'h19d1: q3 = 16'h019a; // 0x33a2
	13'h19d2: q3 = 16'h8701; // 0x33a4
	13'h19d3: q3 = 16'h028a; // 0x33a6
	13'h19d4: q3 = 16'h0666; // 0x33a8
	13'h19d5: q3 = 16'h8a01; // 0x33aa
	13'h19d6: q3 = 16'h019a; // 0x33ac
	13'h19d7: q3 = 16'h8701; // 0x33ae
	13'h19d8: q3 = 16'h0333; // 0x33b0
	13'h19d9: q3 = 16'h0666; // 0x33b2
	13'h19da: q3 = 16'h8a01; // 0x33b4
	13'h19db: q3 = 16'h019a; // 0x33b6
	13'h19dc: q3 = 16'h8701; // 0x33b8
	13'h19dd: q3 = 16'h028a; // 0x33ba
	13'h19de: q3 = 16'h0666; // 0x33bc
	13'h19df: q3 = 16'h8a01; // 0x33be
	13'h19e0: q3 = 16'h019a; // 0x33c0
	13'h19e1: q3 = 16'h8701; // 0x33c2
	13'h19e2: q3 = 16'h0333; // 0x33c4
	13'h19e3: q3 = 16'h0ccc; // 0x33c6
	13'h19e4: q3 = 16'h8a01; // 0x33c8
	13'h19e5: q3 = 16'h0334; // 0x33ca
	13'h19e6: q3 = 16'h8701; // 0x33cc
	13'h19e7: q3 = 16'h0333; // 0x33ce
	13'h19e8: q3 = 16'h0666; // 0x33d0
	13'h19e9: q3 = 16'h8a01; // 0x33d2
	13'h19ea: q3 = 16'h099a; // 0x33d4
	13'h19eb: q3 = 16'h8701; // 0x33d6
	13'h19ec: q3 = 16'h0333; // 0x33d8
	13'h19ed: q3 = 16'h0666; // 0x33da
	13'h19ee: q3 = 16'h8a01; // 0x33dc
	13'h19ef: q3 = 16'h019a; // 0x33de
	13'h19f0: q3 = 16'h8701; // 0x33e0
	13'h19f1: q3 = 16'h0333; // 0x33e2
	13'h19f2: q3 = 16'h0333; // 0x33e4
	13'h19f3: q3 = 16'h8a01; // 0x33e6
	13'h19f4: q3 = 16'h00cd; // 0x33e8
	13'h19f5: q3 = 16'h8701; // 0x33ea
	13'h19f6: q3 = 16'h0333; // 0x33ec
	13'h19f7: q3 = 16'h0333; // 0x33ee
	13'h19f8: q3 = 16'h8a01; // 0x33f0
	13'h19f9: q3 = 16'h00cd; // 0x33f2
	13'h19fa: q3 = 16'h8701; // 0x33f4
	13'h19fb: q3 = 16'h0333; // 0x33f6
	13'h19fc: q3 = 16'h0666; // 0x33f8
	13'h19fd: q3 = 16'h8a01; // 0x33fa
	13'h19fe: q3 = 16'h019a; // 0x33fc
	13'h19ff: q3 = 16'h8701; // 0x33fe
	13'h1a00: q3 = 16'h028a; // 0x3400
	13'h1a01: q3 = 16'h0666; // 0x3402
	13'h1a02: q3 = 16'h8a01; // 0x3404
	13'h1a03: q3 = 16'h019a; // 0x3406
	13'h1a04: q3 = 16'h8701; // 0x3408
	13'h1a05: q3 = 16'h0333; // 0x340a
	13'h1a06: q3 = 16'h0ccc; // 0x340c
	13'h1a07: q3 = 16'h8a01; // 0x340e
	13'h1a08: q3 = 16'h1334; // 0x3410
	13'h1a09: q3 = 16'h0100; // 0x3412
	13'h1a0a: q3 = 16'h8701; // 0x3414
	13'h1a0b: q3 = 16'h028a; // 0x3416
	13'h1a0c: q3 = 16'h0800; // 0x3418
	13'h1a0d: q3 = 16'h8701; // 0x341a
	13'h1a0e: q3 = 16'h0222; // 0x341c
	13'h1a0f: q3 = 16'h0800; // 0x341e
	13'h1a10: q3 = 16'h8701; // 0x3420
	13'h1a11: q3 = 16'h028a; // 0x3422
	13'h1a12: q3 = 16'h0800; // 0x3424
	13'h1a13: q3 = 16'h8701; // 0x3426
	13'h1a14: q3 = 16'h0222; // 0x3428
	13'h1a15: q3 = 16'h0800; // 0x342a
	13'h1a16: q3 = 16'h8701; // 0x342c
	13'h1a17: q3 = 16'h028a; // 0x342e
	13'h1a18: q3 = 16'h1000; // 0x3430
	13'h1a19: q3 = 16'h8701; // 0x3432
	13'h1a1a: q3 = 16'h028a; // 0x3434
	13'h1a1b: q3 = 16'h0800; // 0x3436
	13'h1a1c: q3 = 16'h8a01; // 0x3438
	13'h1a1d: q3 = 16'h0800; // 0x343a
	13'h1a1e: q3 = 16'h8701; // 0x343c
	13'h1a1f: q3 = 16'h028a; // 0x343e
	13'h1a20: q3 = 16'h0800; // 0x3440
	13'h1a21: q3 = 16'h8701; // 0x3442
	13'h1a22: q3 = 16'h028a; // 0x3444
	13'h1a23: q3 = 16'h0400; // 0x3446
	13'h1a24: q3 = 16'h8701; // 0x3448
	13'h1a25: q3 = 16'h028a; // 0x344a
	13'h1a26: q3 = 16'h0400; // 0x344c
	13'h1a27: q3 = 16'h8701; // 0x344e
	13'h1a28: q3 = 16'h028a; // 0x3450
	13'h1a29: q3 = 16'h0800; // 0x3452
	13'h1a2a: q3 = 16'h8701; // 0x3454
	13'h1a2b: q3 = 16'h0222; // 0x3456
	13'h1a2c: q3 = 16'h0800; // 0x3458
	13'h1a2d: q3 = 16'h8701; // 0x345a
	13'h1a2e: q3 = 16'h028a; // 0x345c
	13'h1a2f: q3 = 16'h1000; // 0x345e
	13'h1a30: q3 = 16'h8a01; // 0x3460
	13'h1a31: q3 = 16'h1000; // 0x3462
	13'h1a32: q3 = 16'h8701; // 0x3464
	13'h1a33: q3 = 16'h0445; // 0x3466
	13'h1a34: q3 = 16'h0800; // 0x3468
	13'h1a35: q3 = 16'h8701; // 0x346a
	13'h1a36: q3 = 16'h0333; // 0x346c
	13'h1a37: q3 = 16'h0800; // 0x346e
	13'h1a38: q3 = 16'h8701; // 0x3470
	13'h1a39: q3 = 16'h0445; // 0x3472
	13'h1a3a: q3 = 16'h0800; // 0x3474
	13'h1a3b: q3 = 16'h8701; // 0x3476
	13'h1a3c: q3 = 16'h0333; // 0x3478
	13'h1a3d: q3 = 16'h0800; // 0x347a
	13'h1a3e: q3 = 16'h8701; // 0x347c
	13'h1a3f: q3 = 16'h0445; // 0x347e
	13'h1a40: q3 = 16'h1000; // 0x3480
	13'h1a41: q3 = 16'h8701; // 0x3482
	13'h1a42: q3 = 16'h0445; // 0x3484
	13'h1a43: q3 = 16'h0800; // 0x3486
	13'h1a44: q3 = 16'h8a01; // 0x3488
	13'h1a45: q3 = 16'h0800; // 0x348a
	13'h1a46: q3 = 16'h8701; // 0x348c
	13'h1a47: q3 = 16'h0445; // 0x348e
	13'h1a48: q3 = 16'h0800; // 0x3490
	13'h1a49: q3 = 16'h8701; // 0x3492
	13'h1a4a: q3 = 16'h0445; // 0x3494
	13'h1a4b: q3 = 16'h0400; // 0x3496
	13'h1a4c: q3 = 16'h8701; // 0x3498
	13'h1a4d: q3 = 16'h0445; // 0x349a
	13'h1a4e: q3 = 16'h0400; // 0x349c
	13'h1a4f: q3 = 16'h8701; // 0x349e
	13'h1a50: q3 = 16'h0445; // 0x34a0
	13'h1a51: q3 = 16'h0800; // 0x34a2
	13'h1a52: q3 = 16'h8701; // 0x34a4
	13'h1a53: q3 = 16'h0333; // 0x34a6
	13'h1a54: q3 = 16'h0800; // 0x34a8
	13'h1a55: q3 = 16'h8701; // 0x34aa
	13'h1a56: q3 = 16'h0445; // 0x34ac
	13'h1a57: q3 = 16'h1000; // 0x34ae
	13'h1a58: q3 = 16'h8a01; // 0x34b0
	13'h1a59: q3 = 16'h1000; // 0x34b2
	13'h1a5a: q3 = 16'h0100; // 0x34b4
	13'h1a5b: q3 = 16'h013b; // 0x34b6
	13'h1a5c: q3 = 16'h0195; // 0x34b8
	13'h1a5d: q3 = 16'h01ef; // 0x34ba
	13'h1a5e: q3 = 16'h0249; // 0x34bc
	13'h1a5f: q3 = 16'h02a3; // 0x34be
	13'h1a60: q3 = 16'h02fd; // 0x34c0
	13'h1a61: q3 = 16'h0357; // 0x34c2
	13'h1a62: q3 = 16'h03b1; // 0x34c4
	13'h1a63: q3 = 16'h001b; // 0x34c6
	13'h1a64: q3 = 16'h0023; // 0x34c8
	13'h1a65: q3 = 16'h002b; // 0x34ca
	13'h1a66: q3 = 16'h0037; // 0x34cc
	13'h1a67: q3 = 16'h0043; // 0x34ce
	13'h1a68: q3 = 16'h0049; // 0x34d0
	13'h1a69: q3 = 16'h0053; // 0x34d2
	13'h1a6a: q3 = 16'h005b; // 0x34d4
	13'h1a6b: q3 = 16'h0000; // 0x34d6
	13'h1a6c: q3 = 16'hd0c0; // 0x34d8
	13'h1a6d: q3 = 16'h0000; // 0x34da
	13'h1a6e: q3 = 16'hcf12; // 0x34dc
	13'h1a6f: q3 = 16'h0000; // 0x34de
	13'h1a70: q3 = 16'hcf40; // 0x34e0
	13'h1a71: q3 = 16'h0000; // 0x34e2
	13'h1a72: q3 = 16'hcf74; // 0x34e4
	13'h1a73: q3 = 16'h0000; // 0x34e6
	13'h1a74: q3 = 16'hcfa2; // 0x34e8
	13'h1a75: q3 = 16'h0000; // 0x34ea
	13'h1a76: q3 = 16'hcfee; // 0x34ec
	13'h1a77: q3 = 16'h0000; // 0x34ee
	13'h1a78: q3 = 16'hd02e; // 0x34f0
	13'h1a79: q3 = 16'h0000; // 0x34f2
	13'h1a7a: q3 = 16'hd074; // 0x34f4
	13'h1a7b: q3 = 16'h0000; // 0x34f6
	13'h1a7c: q3 = 16'h7f3a; // 0x34f8
	13'h1a7d: q3 = 16'h0000; // 0x34fa
	13'h1a7e: q3 = 16'h7f5a; // 0x34fc
	13'h1a7f: q3 = 16'h0000; // 0x34fe
	13'h1a80: q3 = 16'h7f78; // 0x3500
	13'h1a81: q3 = 16'h0000; // 0x3502
	13'h1a82: q3 = 16'h7f7a; // 0x3504
	13'h1a83: q3 = 16'h020c; // 0x3506
	13'h1a84: q3 = 16'h161a; // 0x3508
	13'h1a85: q3 = 16'h0610; // 0x350a
	13'h1a86: q3 = 16'h0004; // 0x350c
	13'h1a87: q3 = 16'h0a0e; // 0x350e
	13'h1a88: q3 = 16'h1418; // 0x3510
	13'h1a89: q3 = 16'hff00; // 0x3512
	13'h1a8a: q3 = 16'h000a; // 0x3514
	13'h1a8b: q3 = 16'h1418; // 0x3516
	13'h1a8c: q3 = 16'h0e04; // 0x3518
	13'h1a8d: q3 = 16'hff00; // 0x351a
	13'h1a8e: q3 = 16'h00a4; // 0x351c
	13'h1a8f: q3 = 16'h0000; // 0x351e
	13'h1a90: q3 = 16'h0004; // 0x3520
	13'h1a91: q3 = 16'h0000; // 0x3522
	13'h1a92: q3 = 16'h02d0; // 0x3524
	13'h1a93: q3 = 16'h02d0; // 0x3526
	13'h1a94: q3 = 16'h0010; // 0x3528
	13'h1a95: q3 = 16'h00dc; // 0x352a
	13'h1a96: q3 = 16'h00ce; // 0x352c
	13'h1a97: q3 = 16'h001f; // 0x352e
	13'h1a98: q3 = 16'h0068; // 0x3530
	13'h1a99: q3 = 16'h0057; // 0x3532
	13'h1a9a: q3 = 16'h0029; // 0x3534
	13'h1a9b: q3 = 16'h0000; // 0x3536
	13'h1a9c: q3 = 16'h0000; // 0x3538
	13'h1a9d: q3 = 16'h0000; // 0x353a
	13'h1a9e: q3 = 16'h0780; // 0x353c
	13'h1a9f: q3 = 16'h0780; // 0x353e
	13'h1aa0: q3 = 16'h0001; // 0x3540
	13'h1aa1: q3 = 16'hffe4; // 0x3542
	13'h1aa2: q3 = 16'hffea; // 0x3544
	13'h1aa3: q3 = 16'h0057; // 0x3546
	13'h1aa4: q3 = 16'h0000; // 0x3548
	13'h1aa5: q3 = 16'h02d0; // 0x354a
	13'h1aa6: q3 = 16'h0000; // 0x354c
	13'h1aa7: q3 = 16'h0000; // 0x354e
	13'h1aa8: q3 = 16'h8136; // 0x3550
	13'h1aa9: q3 = 16'h0000; // 0x3552
	13'h1aaa: q3 = 16'hf524; // 0x3554
	13'h1aab: q3 = 16'h2600; // 0x3556
	13'h1aac: q3 = 16'h0000; // 0x3558
	13'h1aad: q3 = 16'h0000; // 0x355a
	13'h1aae: q3 = 16'h8136; // 0x355c
	13'h1aaf: q3 = 16'h0000; // 0x355e
	13'h1ab0: q3 = 16'hf53c; // 0x3560
	13'h1ab1: q3 = 16'h0000; // 0x3562
	13'h1ab2: q3 = 16'h0000; // 0x3564
	13'h1ab3: q3 = 16'h0000; // 0x3566
	13'h1ab4: q3 = 16'h0000; // 0x3568
	13'h1ab5: q3 = 16'h00e0; // 0x356a
	13'h1ab6: q3 = 16'h0000; // 0x356c
	13'h1ab7: q3 = 16'h05d2; // 0x356e
	13'h1ab8: q3 = 16'h0000; // 0x3570
	13'h1ab9: q3 = 16'h0000; // 0x3572
	13'h1aba: q3 = 16'hf54e; // 0x3574
	13'h1abb: q3 = 16'hffff; // 0x3576
	13'h1abc: q3 = 16'hffc6; // 0x3578
	13'h1abd: q3 = 16'hffd5; // 0x357a
	13'h1abe: q3 = 16'h0053; // 0x357c
	13'h1abf: q3 = 16'hff8b; // 0x357e
	13'h1ac0: q3 = 16'hff99; // 0x3580
	13'h1ac1: q3 = 16'h003e; // 0x3582
	13'h1ac2: q3 = 16'hfe7a; // 0x3584
	13'h1ac3: q3 = 16'hfe8d; // 0x3586
	13'h1ac4: q3 = 16'h001f; // 0x3588
	13'h1ac5: q3 = 16'h0000; // 0x358a
	13'h1ac6: q3 = 16'h0000; // 0x358c
	13'h1ac7: q3 = 16'h0000; // 0x358e
	13'h1ac8: q3 = 16'h00b4; // 0x3590
	13'h1ac9: q3 = 16'h000a; // 0x3592
	13'h1aca: q3 = 16'h00af; // 0x3594
	13'h1acb: q3 = 16'hf880; // 0x3596
	13'h1acc: q3 = 16'hf880; // 0x3598
	13'h1acd: q3 = 16'h0001; // 0x359a
	13'h1ace: q3 = 16'h0000; // 0x359c
	13'h1acf: q3 = 16'hffc6; // 0x359e
	13'h1ad0: q3 = 16'h0000; // 0x35a0
	13'h1ad1: q3 = 16'h0000; // 0x35a2
	13'h1ad2: q3 = 16'h8136; // 0x35a4
	13'h1ad3: q3 = 16'h0000; // 0x35a6
	13'h1ad4: q3 = 16'hf578; // 0x35a8
	13'h1ad5: q3 = 16'h7a00; // 0x35aa
	13'h1ad6: q3 = 16'h0000; // 0x35ac
	13'h1ad7: q3 = 16'h0000; // 0x35ae
	13'h1ad8: q3 = 16'h8136; // 0x35b0
	13'h1ad9: q3 = 16'h0000; // 0x35b2
	13'h1ada: q3 = 16'hf590; // 0x35b4
	13'h1adb: q3 = 16'h0000; // 0x35b6
	13'h1adc: q3 = 16'h0000; // 0x35b8
	13'h1add: q3 = 16'h0000; // 0x35ba
	13'h1ade: q3 = 16'h0000; // 0x35bc
	13'h1adf: q3 = 16'h5859; // 0x35be
	13'h1ae0: q3 = 16'h0000; // 0x35c0
	13'h1ae1: q3 = 16'h05dc; // 0x35c2
	13'h1ae2: q3 = 16'h0000; // 0x35c4
	13'h1ae3: q3 = 16'h0000; // 0x35c6
	13'h1ae4: q3 = 16'hf5a2; // 0x35c8
	13'h1ae5: q3 = 16'hffff; // 0x35ca
	13'h1ae6: q3 = 16'h0008; // 0x35cc
	13'h1ae7: q3 = 16'h000e; // 0x35ce
	13'h1ae8: q3 = 16'h0007; // 0x35d0
	13'h1ae9: q3 = 16'h0031; // 0x35d2
	13'h1aea: q3 = 16'h000b; // 0x35d4
	13'h1aeb: q3 = 16'h001c; // 0x35d6
	13'h1aec: q3 = 16'h0015; // 0x35d8
	13'h1aed: q3 = 16'h0004; // 0x35da
	13'h1aee: q3 = 16'h0034; // 0x35dc
	13'h1aef: q3 = 16'hffe6; // 0x35de
	13'h1af0: q3 = 16'h0006; // 0x35e0
	13'h1af1: q3 = 16'h0016; // 0x35e2
	13'h1af2: q3 = 16'h0006; // 0x35e4
	13'h1af3: q3 = 16'h0036; // 0x35e6
	13'h1af4: q3 = 16'h0009; // 0x35e8
	13'h1af5: q3 = 16'h001a; // 0x35ea
	13'h1af6: q3 = 16'h0011; // 0x35ec
	13'h1af7: q3 = 16'h0006; // 0x35ee
	13'h1af8: q3 = 16'h002d; // 0x35f0
	13'h1af9: q3 = 16'hffe8; // 0x35f2
	13'h1afa: q3 = 16'h001b; // 0x35f4
	13'h1afb: q3 = 16'h0008; // 0x35f6
	13'h1afc: q3 = 16'h0001; // 0x35f8
	13'h1afd: q3 = 16'h003c; // 0x35fa
	13'h1afe: q3 = 16'hffe7; // 0x35fc
	13'h1aff: q3 = 16'h0000; // 0x35fe
	13'h1b00: q3 = 16'h0010; // 0x3600
	13'h1b01: q3 = 16'h00ee; // 0x3602
	13'h1b02: q3 = 16'h00a8; // 0x3604
	13'h1b03: q3 = 16'h00a4; // 0x3606
	13'h1b04: q3 = 16'h0027; // 0x3608
	13'h1b05: q3 = 16'hfd40; // 0x360a
	13'h1b06: q3 = 16'hfd40; // 0x360c
	13'h1b07: q3 = 16'h001c; // 0x360e
	13'h1b08: q3 = 16'h0000; // 0x3610
	13'h1b09: q3 = 16'h0000; // 0x3612
	13'h1b0a: q3 = 16'h0000; // 0x3614
	13'h1b0b: q3 = 16'h0034; // 0x3616
	13'h1b0c: q3 = 16'h002e; // 0x3618
	13'h1b0d: q3 = 16'h000b; // 0x361a
	13'h1b0e: q3 = 16'h0000; // 0x361c
	13'h1b0f: q3 = 16'h0000; // 0x361e
	13'h1b10: q3 = 16'h002b; // 0x3620
	13'h1b11: q3 = 16'hffd4; // 0x3622
	13'h1b12: q3 = 16'hffd9; // 0x3624
	13'h1b13: q3 = 16'h000d; // 0x3626
	13'h1b14: q3 = 16'h0000; // 0x3628
	13'h1b15: q3 = 16'h00a8; // 0x362a
	13'h1b16: q3 = 16'h0000; // 0x362c
	13'h1b17: q3 = 16'h0080; // 0x362e
	13'h1b18: q3 = 16'h0050; // 0x3630
	13'h1b19: q3 = 16'h00e0; // 0x3632
	13'h1b1a: q3 = 16'h0000; // 0x3634
	13'h1b1b: q3 = 16'h0000; // 0x3636
	13'h1b1c: q3 = 16'h8136; // 0x3638
	13'h1b1d: q3 = 16'h0000; // 0x363a
	13'h1b1e: q3 = 16'hf604; // 0x363c
	13'h1b1f: q3 = 16'h3400; // 0x363e
	13'h1b20: q3 = 16'h0000; // 0x3640
	13'h1b21: q3 = 16'h0000; // 0x3642
	13'h1b22: q3 = 16'h8136; // 0x3644
	13'h1b23: q3 = 16'h0000; // 0x3646
	13'h1b24: q3 = 16'hf616; // 0x3648
	13'h1b25: q3 = 16'h0000; // 0x364a
	13'h1b26: q3 = 16'h0000; // 0x364c
	13'h1b27: q3 = 16'h0000; // 0x364e
	13'h1b28: q3 = 16'hf62e; // 0x3650
	13'h1b29: q3 = 16'h00e0; // 0x3652
	13'h1b2a: q3 = 16'h0000; // 0x3654
	13'h1b2b: q3 = 16'h00ba; // 0x3656
	13'h1b2c: q3 = 16'h00b1; // 0x3658
	13'h1b2d: q3 = 16'h0027; // 0x365a
	13'h1b2e: q3 = 16'hfebf; // 0x365c
	13'h1b2f: q3 = 16'hfed3; // 0x365e
	13'h1b30: q3 = 16'h001c; // 0x3660
	13'h1b31: q3 = 16'h0000; // 0x3662
	13'h1b32: q3 = 16'h001a; // 0x3664
	13'h1b33: q3 = 16'h0000; // 0x3666
	13'h1b34: q3 = 16'h0070; // 0x3668
	13'h1b35: q3 = 16'h0068; // 0x366a
	13'h1b36: q3 = 16'h000b; // 0x366c
	13'h1b37: q3 = 16'h0000; // 0x366e
	13'h1b38: q3 = 16'h0000; // 0x3670
	13'h1b39: q3 = 16'h0027; // 0x3672
	13'h1b3a: q3 = 16'hffb0; // 0x3674
	13'h1b3b: q3 = 16'hffbd; // 0x3676
	13'h1b3c: q3 = 16'h0011; // 0x3678
	13'h1b3d: q3 = 16'h0000; // 0x367a
	13'h1b3e: q3 = 16'h0080; // 0x367c
	13'h1b3f: q3 = 16'h0000; // 0x367e
	13'h1b40: q3 = 16'h0000; // 0x3680
	13'h1b41: q3 = 16'h8136; // 0x3682
	13'h1b42: q3 = 16'h0000; // 0x3684
	13'h1b43: q3 = 16'hf656; // 0x3686
	13'h1b44: q3 = 16'h0b00; // 0x3688
	13'h1b45: q3 = 16'h0000; // 0x368a
	13'h1b46: q3 = 16'h0000; // 0x368c
	13'h1b47: q3 = 16'h8136; // 0x368e
	13'h1b48: q3 = 16'h0000; // 0x3690
	13'h1b49: q3 = 16'hf668; // 0x3692
	13'h1b4a: q3 = 16'h0000; // 0x3694
	13'h1b4b: q3 = 16'h0000; // 0x3696
	13'h1b4c: q3 = 16'h0000; // 0x3698
	13'h1b4d: q3 = 16'h0000; // 0x369a
	13'h1b4e: q3 = 16'h6c6d; // 0x369c
	13'h1b4f: q3 = 16'h0000; // 0x369e
	13'h1b50: q3 = 16'h0040; // 0x36a0
	13'h1b51: q3 = 16'h005f; // 0x36a2
	13'h1b52: q3 = 16'h0000; // 0x36a4
	13'h1b53: q3 = 16'h0000; // 0x36a6
	13'h1b54: q3 = 16'h0000; // 0x36a8
	13'h1b55: q3 = 16'hf6a0; // 0x36aa
	13'h1b56: q3 = 16'h0000; // 0x36ac
	13'h1b57: q3 = 16'h0000; // 0x36ae
	13'h1b58: q3 = 16'h07c0; // 0x36b0
	13'h1b59: q3 = 16'h0001; // 0x36b2
	13'h1b5a: q3 = 16'h0000; // 0x36b4
	13'h1b5b: q3 = 16'hf636; // 0x36b6
	13'h1b5c: q3 = 16'h0000; // 0x36b8
	13'h1b5d: q3 = 16'hf6a8; // 0x36ba
	13'h1b5e: q3 = 16'h0000; // 0x36bc
	13'h1b5f: q3 = 16'h0000; // 0x36be
	13'h1b60: q3 = 16'hf680; // 0x36c0
	13'h1b61: q3 = 16'hffff; // 0x36c2
	13'h1b62: q3 = 16'h0016; // 0x36c4
	13'h1b63: q3 = 16'h000a; // 0x36c6
	13'h1b64: q3 = 16'h0011; // 0x36c8
	13'h1b65: q3 = 16'h000f; // 0x36ca
	13'h1b66: q3 = 16'h0018; // 0x36cc
	13'h1b67: q3 = 16'h4040; // 0x36ce
	13'h1b68: q3 = 16'h9640; // 0x36d0
	13'h1b69: q3 = 16'h4040; // 0x36d2
	13'h1b6a: q3 = 16'h9696; // 0x36d4
	13'h1b6b: q3 = 16'h4040; // 0x36d6
	13'h1b6c: q3 = 16'h9697; // 0x36d8
	13'h1b6d: q3 = 16'h4040; // 0x36da
	13'h1b6e: q3 = 16'h9797; // 0x36dc
	13'h1b6f: q3 = 16'h9640; // 0x36de
	13'h1b70: q3 = 16'h9797; // 0x36e0
	13'h1b71: q3 = 16'h9696; // 0x36e2
	13'h1b72: q3 = 16'h9797; // 0x36e4
	13'h1b73: q3 = 16'h9697; // 0x36e6
	13'h1b74: q3 = 16'h9797; // 0x36e8
	13'h1b75: q3 = 16'h9797; // 0x36ea
	13'h1b76: q3 = 16'h9797; // 0x36ec
	13'h1b77: q3 = 16'h4040; // 0x36ee
	13'h1b78: q3 = 16'h9040; // 0x36f0
	13'h1b79: q3 = 16'h4040; // 0x36f2
	13'h1b7a: q3 = 16'h9090; // 0x36f4
	13'h1b7b: q3 = 16'h4040; // 0x36f6
	13'h1b7c: q3 = 16'h9091; // 0x36f8
	13'h1b7d: q3 = 16'h4040; // 0x36fa
	13'h1b7e: q3 = 16'h9191; // 0x36fc
	13'h1b7f: q3 = 16'h9040; // 0x36fe
	13'h1b80: q3 = 16'h9191; // 0x3700
	13'h1b81: q3 = 16'h9090; // 0x3702
	13'h1b82: q3 = 16'h9191; // 0x3704
	13'h1b83: q3 = 16'h9091; // 0x3706
	13'h1b84: q3 = 16'h9191; // 0x3708
	13'h1b85: q3 = 16'h9191; // 0x370a
	13'h1b86: q3 = 16'h9191; // 0x370c
	13'h1b87: q3 = 16'hb8b9; // 0x370e
	13'h1b88: q3 = 16'hbabb; // 0x3710
	13'h1b89: q3 = 16'hbcbd; // 0x3712
	13'h1b8a: q3 = 16'hbebf; // 0x3714
	13'h1b8b: q3 = 16'hc0c1; // 0x3716
	13'h1b8c: q3 = 16'hc2c3; // 0x3718
	13'h1b8d: q3 = 16'hc4c5; // 0x371a
	13'h1b8e: q3 = 16'hc6c7; // 0x371c
	13'h1b8f: q3 = 16'hc8c9; // 0x371e
	13'h1b90: q3 = 16'hcacb; // 0x3720
	13'h1b91: q3 = 16'hcccd; // 0x3722
	13'h1b92: q3 = 16'hcecf; // 0x3724
	13'h1b93: q3 = 16'hd0d1; // 0x3726
	13'h1b94: q3 = 16'hd2d3; // 0x3728
	13'h1b95: q3 = 16'hd4d5; // 0x372a
	13'h1b96: q3 = 16'hd6d7; // 0x372c
	13'h1b97: q3 = 16'h9899; // 0x372e
	13'h1b98: q3 = 16'h9a9b; // 0x3730
	13'h1b99: q3 = 16'h9c9d; // 0x3732
	13'h1b9a: q3 = 16'h9e9f; // 0x3734
	13'h1b9b: q3 = 16'ha0a1; // 0x3736
	13'h1b9c: q3 = 16'ha2a3; // 0x3738
	13'h1b9d: q3 = 16'ha4a5; // 0x373a
	13'h1b9e: q3 = 16'ha6a7; // 0x373c
	13'h1b9f: q3 = 16'ha8a9; // 0x373e
	13'h1ba0: q3 = 16'haaab; // 0x3740
	13'h1ba1: q3 = 16'hacad; // 0x3742
	13'h1ba2: q3 = 16'haeaf; // 0x3744
	13'h1ba3: q3 = 16'hb0b1; // 0x3746
	13'h1ba4: q3 = 16'hb2b3; // 0x3748
	13'h1ba5: q3 = 16'hb4b5; // 0x374a
	13'h1ba6: q3 = 16'hb6b7; // 0x374c
	13'h1ba7: q3 = 16'h1011; // 0x374e
	13'h1ba8: q3 = 16'h1213; // 0x3750
	13'h1ba9: q3 = 16'h1011; // 0x3752
	13'h1baa: q3 = 16'h1213; // 0x3754
	13'h1bab: q3 = 16'h1011; // 0x3756
	13'h1bac: q3 = 16'h1213; // 0x3758
	13'h1bad: q3 = 16'h1011; // 0x375a
	13'h1bae: q3 = 16'h1213; // 0x375c
	13'h1baf: q3 = 16'h1011; // 0x375e
	13'h1bb0: q3 = 16'h1213; // 0x3760
	13'h1bb1: q3 = 16'h1011; // 0x3762
	13'h1bb2: q3 = 16'h1213; // 0x3764
	13'h1bb3: q3 = 16'h1011; // 0x3766
	13'h1bb4: q3 = 16'h1213; // 0x3768
	13'h1bb5: q3 = 16'h1011; // 0x376a
	13'h1bb6: q3 = 16'h1213; // 0x376c
	13'h1bb7: q3 = 16'h2020; // 0x376e
	13'h1bb8: q3 = 16'h3000; // 0x3770
	13'h1bb9: q3 = 16'h3000; // 0x3772
	13'h1bba: q3 = 16'h0000; // 0x3774
	13'h1bbb: q3 = 16'h0078; // 0x3776
	13'h1bbc: q3 = 16'h0000; // 0x3778
	13'h1bbd: q3 = 16'h00a8; // 0x377a
	13'h1bbe: q3 = 16'h0000; // 0x377c
	13'h1bbf: q3 = 16'h0a12; // 0x377e
	13'h1bc0: q3 = 16'h0f11; // 0x3780
	13'h1bc1: q3 = 16'h280b; // 0x3782
	13'h1bc2: q3 = 16'h1f64; // 0x3784
	13'h1bc3: q3 = 16'h0032; // 0x3786
	13'h1bc4: q3 = 16'h0c1e; // 0x3788
	13'h1bc5: q3 = 16'h6400; // 0x378a
	13'h1bc6: q3 = 16'h310d; // 0x378c
	13'h1bc7: q3 = 16'h1d64; // 0x378e
	13'h1bc8: q3 = 16'h0033; // 0x3790
	13'h1bc9: q3 = 16'h0f07; // 0x3792
	13'h1bca: q3 = 16'h6420; // 0x3794
	13'h1bcb: q3 = 16'h3217; // 0x3796
	13'h1bcc: q3 = 16'h1802; // 0x3798
	13'h1bcd: q3 = 16'h003e; // 0x379a
	13'h1bce: q3 = 16'h1a07; // 0x379c
	13'h1bcf: q3 = 16'h6420; // 0x379e
	13'h1bd0: q3 = 16'h321b; // 0x37a0
	13'h1bd1: q3 = 16'h0664; // 0x37a2
	13'h1bd2: q3 = 16'h2032; // 0x37a4
	13'h1bd3: q3 = 16'h1c05; // 0x37a6
	13'h1bd4: q3 = 16'h6420; // 0x37a8
	13'h1bd5: q3 = 16'h2e1d; // 0x37aa
	13'h1bd6: q3 = 16'h0464; // 0x37ac
	13'h1bd7: q3 = 16'h2033; // 0x37ae
	13'h1bd8: q3 = 16'h1e07; // 0x37b0
	13'h1bd9: q3 = 16'h6420; // 0x37b2
	13'h1bda: q3 = 16'h381f; // 0x37b4
	13'h1bdb: q3 = 16'h0664; // 0x37b6
	13'h1bdc: q3 = 16'h2038; // 0x37b8
	13'h1bdd: q3 = 16'h2005; // 0x37ba
	13'h1bde: q3 = 16'h6420; // 0x37bc
	13'h1bdf: q3 = 16'h3121; // 0x37be
	13'h1be0: q3 = 16'h0664; // 0x37c0
	13'h1be1: q3 = 16'h203a; // 0x37c2
	13'h1be2: q3 = 16'h2205; // 0x37c4
	13'h1be3: q3 = 16'h6420; // 0x37c6
	13'h1be4: q3 = 16'h3a23; // 0x37c8
	13'h1be5: q3 = 16'h0664; // 0x37ca
	13'h1be6: q3 = 16'h203c; // 0x37cc
	13'h1be7: q3 = 16'h2405; // 0x37ce
	13'h1be8: q3 = 16'h6420; // 0x37d0
	13'h1be9: q3 = 16'h3c25; // 0x37d2
	13'h1bea: q3 = 16'h0764; // 0x37d4
	13'h1beb: q3 = 16'h2038; // 0x37d6
	13'h1bec: q3 = 16'h2606; // 0x37d8
	13'h1bed: q3 = 16'h6420; // 0x37da
	13'h1bee: q3 = 16'h3127; // 0x37dc
	13'h1bef: q3 = 16'h0764; // 0x37de
	13'h1bf0: q3 = 16'h203c; // 0x37e0
	13'h1bf1: q3 = 16'h2806; // 0x37e2
	13'h1bf2: q3 = 16'h6420; // 0x37e4
	13'h1bf3: q3 = 16'h3c18; // 0x37e6
	13'h1bf4: q3 = 16'h0902; // 0x37e8
	13'h1bf5: q3 = 16'h0031; // 0x37ea
	13'h1bf6: q3 = 16'h1906; // 0x37ec
	13'h1bf7: q3 = 16'h6420; // 0x37ee
	13'h1bf8: q3 = 16'h3c31; // 0x37f0
	13'h1bf9: q3 = 16'h0564; // 0x37f2
	13'h1bfa: q3 = 16'h0031; // 0x37f4
	13'h1bfb: q3 = 16'h3204; // 0x37f6
	13'h1bfc: q3 = 16'h6400; // 0x37f8
	13'h1bfd: q3 = 16'h3134; // 0x37fa
	13'h1bfe: q3 = 16'h1264; // 0x37fc
	13'h1bff: q3 = 16'h0031; // 0x37fe
	13'h1c00: q3 = 16'h3612; // 0x3800
	13'h1c01: q3 = 16'h6400; // 0x3802
	13'h1c02: q3 = 16'h310a; // 0x3804
	13'h1c03: q3 = 16'h0400; // 0x3806
	13'h1c04: q3 = 16'h0028; // 0x3808
	13'h1c05: q3 = 16'h2831; // 0x380a
	13'h1c06: q3 = 16'h2920; // 0x380c
	13'h1c07: q3 = 16'h0028; // 0x380e
	13'h1c08: q3 = 16'h3229; // 0x3810
	13'h1c09: q3 = 16'h2000; // 0x3812
	13'h1c0a: q3 = 16'h2000; // 0x3814
	13'h1c0b: q3 = 16'h0000; // 0x3816
	13'h1c0c: q3 = 16'h0014; // 0x3818
	13'h1c0d: q3 = 16'h0000; // 0x381a
	13'h1c0e: q3 = 16'h001e; // 0x381c
	13'h1c0f: q3 = 16'h0000; // 0x381e
	13'h1c10: q3 = 16'h0007; // 0x3820
	13'h1c11: q3 = 16'h0767; // 0x3822
	13'h1c12: q3 = 16'h070e; // 0x3824
	13'h1c13: q3 = 16'h0c5f; // 0x3826
	13'h1c14: q3 = 16'h5e55; // 0x3828
	13'h1c15: q3 = 16'h2021; // 0x382a
	13'h1c16: q3 = 16'h18ff; // 0x382c
	13'h1c17: q3 = 16'h9b67; // 0x382e
	13'h1c18: q3 = 16'h3f37; // 0x3830
	13'h1c19: q3 = 16'h2eff; // 0x3832
	13'h1c1a: q3 = 16'hc067; // 0x3834
	13'h1c1b: q3 = 16'hff6f; // 0x3836
	13'h1c1c: q3 = 16'h52ff; // 0x3838
	13'h1c1d: q3 = 16'hfead; // 0x383a
	13'h1c1e: q3 = 16'hffae; // 0x383c
	13'h1c1f: q3 = 16'h14ff; // 0x383e
	13'h1c20: q3 = 16'h2818; // 0x3840
	13'h1c21: q3 = 16'h1414; // 0x3842
	13'h1c22: q3 = 16'h0b2e; // 0x3844
	13'h1c23: q3 = 16'h3f67; // 0x3846
	13'h1c24: q3 = 16'hff07; // 0x3848
	13'h1c25: q3 = 16'h0417; // 0x384a
	13'h1c26: q3 = 16'h156f; // 0x384c
	13'h1c27: q3 = 16'hff5f; // 0x384e
	13'h1c28: q3 = 16'h5220; // 0x3850
	13'h1c29: q3 = 16'h2010; // 0x3852
	13'h1c2a: q3 = 16'hff13; // 0x3854
	13'h1c2b: q3 = 16'h0a3f; // 0x3856
	13'h1c2c: q3 = 16'h3f67; // 0x3858
	13'h1c2d: q3 = 16'hff4e; // 0x385a
	13'h1c2e: q3 = 16'h5490; // 0x385c
	13'h1c2f: q3 = 16'he067; // 0x385e
	13'h1c30: q3 = 16'h3f27; // 0x3860
	13'h1c31: q3 = 16'h1552; // 0x3862
	13'h1c32: q3 = 16'h5252; // 0x3864
	13'h1c33: q3 = 16'h077a; // 0x3866
	13'h1c34: q3 = 16'h52ff; // 0x3868
	13'h1c35: q3 = 16'h3f26; // 0x386a
	13'h1c36: q3 = 16'h1414; // 0x386c
	13'h1c37: q3 = 16'h6720; // 0x386e
	13'h1c38: q3 = 16'h2067; // 0x3870
	13'h1c39: q3 = 16'h5f5f; // 0x3872
	13'h1c3a: q3 = 16'h672e; // 0x3874
	13'h1c3b: q3 = 16'h3f15; // 0x3876
	13'h1c3c: q3 = 16'h0407; // 0x3878
	13'h1c3d: q3 = 16'h67ff; // 0x387a
	13'h1c3e: q3 = 16'had5b; // 0x387c
	13'h1c3f: q3 = 16'ha7a7; // 0x387e
	13'h1c40: q3 = 16'ha7ff; // 0x3880
	13'h1c41: q3 = 16'h131d; // 0x3882
	13'h1c42: q3 = 16'h6666; // 0x3884
	13'h1c43: q3 = 16'h66b9; // 0x3886
	13'h1c44: q3 = 16'hb9b9; // 0x3888
	13'h1c45: q3 = 16'h8e8e; // 0x388a
	13'h1c46: q3 = 16'h8e51; // 0x388c
	13'h1c47: q3 = 16'h9bff; // 0x388e
	13'h1c48: q3 = 16'h0204; // 0x3890
	13'h1c49: q3 = 16'h0741; // 0x3892
	13'h1c4a: q3 = 16'h4952; // 0x3894
	13'h1c4b: q3 = 16'h121c; // 0x3896
	13'h1c4c: q3 = 16'h2f10; // 0x3898
	13'h1c4d: q3 = 16'h1820; // 0x389a
	13'h1c4e: q3 = 16'h0049; // 0x389c
	13'h1c4f: q3 = 16'h522e; // 0x389e
	13'h1c50: q3 = 16'h3f67; // 0x38a0
	13'h1c51: q3 = 16'h1b2d; // 0x38a2
	13'h1c52: q3 = 16'h3f02; // 0x38a4
	13'h1c53: q3 = 16'h0407; // 0x38a6
	13'h1c54: q3 = 16'h1364; // 0x38a8
	13'h1c55: q3 = 16'h6f41; // 0x38aa
	13'h1c56: q3 = 16'h54a7; // 0x38ac
	13'h1c57: q3 = 16'h0a14; // 0x38ae
	13'h1c58: q3 = 16'h1f12; // 0x38b0
	13'h1c59: q3 = 16'h263f; // 0x38b2
	13'h1c5a: q3 = 16'h121c; // 0x38b4
	13'h1c5b: q3 = 16'h2f0a; // 0x38b6
	13'h1c5c: q3 = 16'h1427; // 0x38b8
	13'h1c5d: q3 = 16'h020b; // 0x38ba
	13'h1c5e: q3 = 16'h1448; // 0x38bc
	13'h1c5f: q3 = 16'h5a6a; // 0x38be
	13'h1c60: q3 = 16'h1020; // 0x38c0
	13'h1c61: q3 = 16'h3858; // 0x38c2
	13'h1c62: q3 = 16'h617a; // 0x38c4
	13'h1c63: q3 = 16'h1018; // 0x38c6
	13'h1c64: q3 = 16'h2040; // 0x38c8
	13'h1c65: q3 = 16'h80c0; // 0x38ca
	13'h1c66: q3 = 16'h8aa0; // 0x38cc
	13'h1c67: q3 = 16'hf040; // 0x38ce
	13'h1c68: q3 = 16'h5180; // 0x38d0
	13'h1c69: q3 = 16'h424d; // 0x38d2
	13'h1c6a: q3 = 16'h4f49; // 0x38d4
	13'h1c6b: q3 = 16'h93c6; // 0x38d6
	13'h1c6c: q3 = 16'h52ac; // 0x38d8
	13'h1c6d: q3 = 16'hff48; // 0x38da
	13'h1c6e: q3 = 16'h4952; // 0x38dc
	13'h1c6f: q3 = 16'h05f5; // 0x38de
	13'h1c70: q3 = 16'he0ff; // 0x38e0
	13'h1c71: q3 = 16'h05f5; // 0x38e2
	13'h1c72: q3 = 16'he100; // 0x38e4
	13'h1c73: q3 = 16'h3030; // 0x38e6
	13'h1c74: q3 = 16'h0030; // 0x38e8
	13'h1c75: q3 = 16'h3000; // 0x38ea
	13'h1c76: q3 = 16'h0000; // 0x38ec
	13'h1c77: q3 = 16'h003c; // 0x38ee
	13'h1c78: q3 = 16'h4a41; // 0x38f0
	13'h1c79: q3 = 16'h4854; // 0x38f2
	13'h1c7a: q3 = 16'h5720; // 0x38f4
	13'h1c7b: q3 = 16'h5242; // 0x38f6
	13'h1c7c: q3 = 16'h4a4a; // 0x38f8
	13'h1c7d: q3 = 16'h4148; // 0x38fa
	13'h1c7e: q3 = 16'h5457; // 0x38fc
	13'h1c7f: q3 = 16'h2052; // 0x38fe
	13'h1c80: q3 = 16'h424a; // 0x3900
	13'h1c81: q3 = 16'h4247; // 0x3902
	13'h1c82: q3 = 16'h424c; // 0x3904
	13'h1c83: q3 = 16'h5244; // 0x3906
	13'h1c84: q3 = 16'h5052; // 0x3908
	13'h1c85: q3 = 16'h4752; // 0x390a
	13'h1c86: q3 = 16'h4f59; // 0x390c
	13'h1c87: q3 = 16'h4445; // 0x390e
	13'h1c88: q3 = 16'h4c44; // 0x3910
	13'h1c89: q3 = 16'h4f47; // 0x3912
	13'h1c8a: q3 = 16'h4159; // 0x3914
	13'h1c8b: q3 = 16'h4e45; // 0x3916
	13'h1c8c: q3 = 16'h4456; // 0x3918
	13'h1c8d: q3 = 16'h4d4f; // 0x391a
	13'h1c8e: q3 = 16'h4500; // 0x391c
	13'h1c8f: q3 = 16'h021a; // 0x391e
	13'h1c90: q3 = 16'h01dc; // 0x3920
	13'h1c91: q3 = 16'h0194; // 0x3922
	13'h1c92: q3 = 16'h017e; // 0x3924
	13'h1c93: q3 = 16'h0176; // 0x3926
	13'h1c94: q3 = 16'h0171; // 0x3928
	13'h1c95: q3 = 16'h0157; // 0x392a
	13'h1c96: q3 = 16'h0155; // 0x392c
	13'h1c97: q3 = 16'h0153; // 0x392e
	13'h1c98: q3 = 16'h0151; // 0x3930
	13'h1c99: q3 = 16'h013e; // 0x3932
	13'h1c9a: q3 = 16'h013c; // 0x3934
	13'h1c9b: q3 = 16'h0137; // 0x3936
	13'h1c9c: q3 = 16'h0134; // 0x3938
	13'h1c9d: q3 = 16'h012f; // 0x393a
	13'h1c9e: q3 = 16'h0f0e; // 0x393c
	13'h1c9f: q3 = 16'h0d0c; // 0x393e
	13'h1ca0: q3 = 16'h0b0a; // 0x3940
	13'h1ca1: q3 = 16'h0908; // 0x3942
	13'h1ca2: q3 = 16'h0706; // 0x3944
	13'h1ca3: q3 = 16'h0504; // 0x3946
	13'h1ca4: q3 = 16'h0302; // 0x3948
	13'h1ca5: q3 = 16'h0100; // 0x394a
	13'h1ca6: q3 = 16'h0000; // 0x394c
	13'h1ca7: q3 = 16'h000a; // 0x394e
	13'h1ca8: q3 = 16'h0014; // 0x3950
	13'h1ca9: q3 = 16'h001e; // 0x3952
	13'h1caa: q3 = 16'h0028; // 0x3954
	13'h1cab: q3 = 16'h0032; // 0x3956
	13'h1cac: q3 = 16'h003c; // 0x3958
	13'h1cad: q3 = 16'h0046; // 0x395a
	13'h1cae: q3 = 16'h0050; // 0x395c
	13'h1caf: q3 = 16'h005a; // 0x395e
	13'h1cb0: q3 = 16'h0064; // 0x3960
	13'h1cb1: q3 = 16'h006e; // 0x3962
	13'h1cb2: q3 = 16'h0078; // 0x3964
	13'h1cb3: q3 = 16'h007d; // 0x3966
	13'h1cb4: q3 = 16'h03e7; // 0x3968
	13'h1cb5: q3 = 16'h0000; // 0x396a
	13'h1cb6: q3 = 16'h0010; // 0x396c
	13'h1cb7: q3 = 16'h0080; // 0x396e
	13'h1cb8: q3 = 16'h0002; // 0x3970
	13'h1cb9: q3 = 16'h001f; // 0x3972
	13'h1cba: q3 = 16'ha28e; // 0x3974
	13'h1cbb: q3 = 16'h0000; // 0x3976
	13'h1cbc: q3 = 16'h8120; // 0x3978
	13'h1cbd: q3 = 16'h2000; // 0x397a
	13'h1cbe: q3 = 16'h191a; // 0x397c
	13'h1cbf: q3 = 16'h1b1c; // 0x397e
	13'h1cc0: q3 = 16'h1d1e; // 0x3980
	13'h1cc1: q3 = 16'h1fee; // 0x3982
	13'h1cc2: q3 = 16'hecec; // 0x3984
	13'h1cc3: q3 = 16'hecec; // 0x3986
	13'h1cc4: q3 = 16'hecf0; // 0x3988
	13'h1cc5: q3 = 16'h20ed; // 0x398a
	13'h1cc6: q3 = 16'hecec; // 0x398c
	13'h1cc7: q3 = 16'hecef; // 0x398e
	13'h1cc8: q3 = 16'h2020; // 0x3990
	13'h1cc9: q3 = 16'heeec; // 0x3992
	13'h1cca: q3 = 16'hecec; // 0x3994
	13'h1ccb: q3 = 16'hf020; // 0x3996
	13'h1ccc: q3 = 16'h2020; // 0x3998
	13'h1ccd: q3 = 16'hedec; // 0x399a
	13'h1cce: q3 = 16'hef20; // 0x399c
	13'h1ccf: q3 = 16'h2020; // 0x399e
	13'h1cd0: q3 = 16'h20ee; // 0x39a0
	13'h1cd1: q3 = 16'hecf0; // 0x39a2
	13'h1cd2: q3 = 16'h2020; // 0x39a4
	13'h1cd3: q3 = 16'h2020; // 0x39a6
	13'h1cd4: q3 = 16'h20f4; // 0x39a8
	13'h1cd5: q3 = 16'h2020; // 0x39aa
	13'h1cd6: q3 = 16'h2000; // 0x39ac
	13'h1cd7: q3 = 16'h0059; // 0x39ae
	13'h1cd8: q3 = 16'h0014; // 0x39b0
	13'h1cd9: q3 = 16'h0012; // 0x39b2
	13'h1cda: q3 = 16'h0010; // 0x39b4
	13'h1cdb: q3 = 16'h001c; // 0x39b6
	13'h1cdc: q3 = 16'h0019; // 0x39b8
	13'h1cdd: q3 = 16'h0017; // 0x39ba
	13'h1cde: q3 = 16'h000d; // 0x39bc
	13'h1cdf: q3 = 16'h0060; // 0x39be
	13'h1ce0: q3 = 16'h0014; // 0x39c0
	13'h1ce1: q3 = 16'h0012; // 0x39c2
	13'h1ce2: q3 = 16'h0010; // 0x39c4
	13'h1ce3: q3 = 16'h000e; // 0x39c6
	13'h1ce4: q3 = 16'h000c; // 0x39c8
	13'h1ce5: q3 = 16'h0019; // 0x39ca
	13'h1ce6: q3 = 16'h0017; // 0x39cc
	13'h1ce7: q3 = 16'h0067; // 0x39ce
	13'h1ce8: q3 = 16'h0019; // 0x39d0
	13'h1ce9: q3 = 16'h0016; // 0x39d2
	13'h1cea: q3 = 16'h0014; // 0x39d4
	13'h1ceb: q3 = 16'h0011; // 0x39d6
	13'h1cec: q3 = 16'h0010; // 0x39d8
	13'h1ced: q3 = 16'h000e; // 0x39da
	13'h1cee: q3 = 16'h006d; // 0x39dc
	13'h1cef: q3 = 16'h0019; // 0x39de
	13'h1cf0: q3 = 16'h0014; // 0x39e0
	13'h1cf1: q3 = 16'h000e; // 0x39e2
	13'h1cf2: q3 = 16'h0070; // 0x39e4
	13'h1cf3: q3 = 16'h001d; // 0x39e6
	13'h1cf4: q3 = 16'h001b; // 0x39e8
	13'h1cf5: q3 = 16'h0018; // 0x39ea
	13'h1cf6: q3 = 16'h0016; // 0x39ec
	13'h1cf7: q3 = 16'h0014; // 0x39ee
	13'h1cf8: q3 = 16'h0012; // 0x39f0
	13'h1cf9: q3 = 16'h0011; // 0x39f2
	13'h1cfa: q3 = 16'h0010; // 0x39f4
	13'h1cfb: q3 = 16'h000e; // 0x39f6
	13'h1cfc: q3 = 16'h000c; // 0x39f8
	13'h1cfd: q3 = 16'h000a; // 0x39fa
	13'h1cfe: q3 = 16'h0007; // 0x39fc
	13'h1cff: q3 = 16'h0014; // 0x39fe
	13'h1d00: q3 = 16'h0012; // 0x3a00
	13'h1d01: q3 = 16'h0011; // 0x3a02
	13'h1d02: q3 = 16'h0010; // 0x3a04
	13'h1d03: q3 = 16'h0000; // 0x3a06
	13'h1d04: q3 = 16'h9d58; // 0x3a08
	13'h1d05: q3 = 16'h0000; // 0x3a0a
	13'h1d06: q3 = 16'h9d60; // 0x3a0c
	13'h1d07: q3 = 16'h0000; // 0x3a0e
	13'h1d08: q3 = 16'h9d68; // 0x3a10
	13'h1d09: q3 = 16'h0080; // 0x3a12
	13'h1d0a: q3 = 16'h001f; // 0x3a14
	13'h1d0b: q3 = 16'h001d; // 0x3a16
	13'h1d0c: q3 = 16'h001b; // 0x3a18
	13'h1d0d: q3 = 16'h0019; // 0x3a1a
	13'h1d0e: q3 = 16'h0017; // 0x3a1c
	13'h1d0f: q3 = 16'h000b; // 0x3a1e
	13'h1d10: q3 = 16'h0007; // 0x3a20
	13'h1d11: q3 = 16'h0087; // 0x3a22
	13'h1d12: q3 = 16'h0016; // 0x3a24
	13'h1d13: q3 = 16'h0015; // 0x3a26
	13'h1d14: q3 = 16'h0014; // 0x3a28
	13'h1d15: q3 = 16'h0013; // 0x3a2a
	13'h1d16: q3 = 16'h0012; // 0x3a2c
	13'h1d17: q3 = 16'h0011; // 0x3a2e
	13'h1d18: q3 = 16'h0010; // 0x3a30
	13'h1d19: q3 = 16'h000f; // 0x3a32
	13'h1d1a: q3 = 16'h000e; // 0x3a34
	13'h1d1b: q3 = 16'h000d; // 0x3a36
	13'h1d1c: q3 = 16'h000a; // 0x3a38
	13'h1d1d: q3 = 16'h0009; // 0x3a3a
	13'h1d1e: q3 = 16'h0006; // 0x3a3c
	13'h1d1f: q3 = 16'h0005; // 0x3a3e
	13'h1d20: q3 = 16'h0004; // 0x3a40
	13'h1d21: q3 = 16'h0005; // 0x3a42
	13'h1d22: q3 = 16'h00c9; // 0x3a44
	13'h1d23: q3 = 16'h00c9; // 0x3a46
	13'h1d24: q3 = 16'h0002; // 0x3a48
	13'h1d25: q3 = 16'h0004; // 0x3a4a
	13'h1d26: q3 = 16'h0002; // 0x3a4c
	13'h1d27: q3 = 16'h0004; // 0x3a4e
	13'h1d28: q3 = 16'h0002; // 0x3a50
	13'h1d29: q3 = 16'h0002; // 0x3a52
	13'h1d2a: q3 = 16'h0003; // 0x3a54
	13'h1d2b: q3 = 16'h0003; // 0x3a56
	13'h1d2c: q3 = 16'h0003; // 0x3a58
	13'h1d2d: q3 = 16'h0003; // 0x3a5a
	13'h1d2e: q3 = 16'h0001; // 0x3a5c
	13'h1d2f: q3 = 16'h0000; // 0x3a5e
	13'h1d30: q3 = 16'h0000; // 0x3a60
	13'h1d31: q3 = 16'h0000; // 0x3a62
	13'h1d32: q3 = 16'h0005; // 0x3a64
	13'h1d33: q3 = 16'h0007; // 0x3a66
	13'h1d34: q3 = 16'h0005; // 0x3a68
	13'h1d35: q3 = 16'h000b; // 0x3a6a
	13'h1d36: q3 = 16'h0005; // 0x3a6c
	13'h1d37: q3 = 16'h000f; // 0x3a6e
	13'h1d38: q3 = 16'h0011; // 0x3a70
	13'h1d39: q3 = 16'h0011; // 0x3a72
	13'h1d3a: q3 = 16'h0014; // 0x3a74
	13'h1d3b: q3 = 16'h0014; // 0x3a76
	13'h1d3c: q3 = 16'h0095; // 0x3a78
	13'h1d3d: q3 = 16'h3030; // 0x3a7a
	13'h1d3e: q3 = 16'h004f; // 0x3a7c
	13'h1d3f: q3 = 16'h4646; // 0x3a7e
	13'h1d40: q3 = 16'h0000; // 0x3a80
	13'h1d41: q3 = 16'h0094; // 0x3a82
	13'h1d42: q3 = 16'h8000; // 0x3a84
	13'h1d43: q3 = 16'h0000; // 0x3a86
	13'h1d44: q3 = 16'ha328; // 0x3a88
	13'h1d45: q3 = 16'h0000; // 0x3a8a
	13'h1d46: q3 = 16'ha33a; // 0x3a8c
	13'h1d47: q3 = 16'h0000; // 0x3a8e
	13'h1d48: q3 = 16'ha34c; // 0x3a90
	13'h1d49: q3 = 16'h0000; // 0x3a92
	13'h1d4a: q3 = 16'ha3dc; // 0x3a94
	13'h1d4b: q3 = 16'h0000; // 0x3a96
	13'h1d4c: q3 = 16'ha35e; // 0x3a98
	13'h1d4d: q3 = 16'h0000; // 0x3a9a
	13'h1d4e: q3 = 16'ha368; // 0x3a9c
	13'h1d4f: q3 = 16'h0000; // 0x3a9e
	13'h1d50: q3 = 16'ha372; // 0x3aa0
	13'h1d51: q3 = 16'h0000; // 0x3aa2
	13'h1d52: q3 = 16'ha382; // 0x3aa4
	13'h1d53: q3 = 16'h0000; // 0x3aa6
	13'h1d54: q3 = 16'ha392; // 0x3aa8
	13'h1d55: q3 = 16'h0000; // 0x3aaa
	13'h1d56: q3 = 16'ha3a2; // 0x3aac
	13'h1d57: q3 = 16'h0000; // 0x3aae
	13'h1d58: q3 = 16'ha3a4; // 0x3ab0
	13'h1d59: q3 = 16'h0000; // 0x3ab2
	13'h1d5a: q3 = 16'ha3dc; // 0x3ab4
	13'h1d5b: q3 = 16'h0000; // 0x3ab6
	13'h1d5c: q3 = 16'ha3b4; // 0x3ab8
	13'h1d5d: q3 = 16'h0000; // 0x3aba
	13'h1d5e: q3 = 16'ha3bc; // 0x3abc
	13'h1d5f: q3 = 16'h0000; // 0x3abe
	13'h1d60: q3 = 16'ha584; // 0x3ac0
	13'h1d61: q3 = 16'h0000; // 0x3ac2
	13'h1d62: q3 = 16'ha58c; // 0x3ac4
	13'h1d63: q3 = 16'h0000; // 0x3ac6
	13'h1d64: q3 = 16'ha594; // 0x3ac8
	13'h1d65: q3 = 16'h0000; // 0x3aca
	13'h1d66: q3 = 16'ha59c; // 0x3acc
	13'h1d67: q3 = 16'h0000; // 0x3ace
	13'h1d68: q3 = 16'ha5a4; // 0x3ad0
	13'h1d69: q3 = 16'h0016; // 0x3ad2
	13'h1d6a: q3 = 16'h2c42; // 0x3ad4
	13'h1d6b: q3 = 16'h586c; // 0x3ad6
	13'h1d6c: q3 = 16'h8093; // 0x3ad8
	13'h1d6d: q3 = 16'ha5b5; // 0x3ada
	13'h1d6e: q3 = 16'hc4d2; // 0x3adc
	13'h1d6f: q3 = 16'hdee8; // 0x3ade
	13'h1d70: q3 = 16'hf1f7; // 0x3ae0
	13'h1d71: q3 = 16'hfcff; // 0x3ae2
	13'h1d72: q3 = 16'h00ff; // 0x3ae4
	13'h1d73: q3 = 16'hfcf7; // 0x3ae6
	13'h1d74: q3 = 16'hf1e8; // 0x3ae8
	13'h1d75: q3 = 16'hded2; // 0x3aea
	13'h1d76: q3 = 16'hc4b5; // 0x3aec
	13'h1d77: q3 = 16'ha593; // 0x3aee
	13'h1d78: q3 = 16'h806c; // 0x3af0
	13'h1d79: q3 = 16'h5842; // 0x3af2
	13'h1d7a: q3 = 16'h2c16; // 0x3af4
	13'h1d7b: q3 = 16'h0d00; // 0x3af6
	13'h1d7c: q3 = 16'h0000; // 0x3af8
	13'h1d7d: q3 = 16'hf386; // 0x3afa
	13'h1d7e: q3 = 16'h0801; // 0x3afc
	13'h1d7f: q3 = 16'h0100; // 0x3afe
	13'h1d80: q3 = 16'h0000; // 0x3b00
	13'h1d81: q3 = 16'h0000; // 0x3b02
	13'h1d82: q3 = 16'h0000; // 0x3b04
	13'h1d83: q3 = 16'hffa8; // 0x3b06
	13'h1d84: q3 = 16'hffb2; // 0x3b08
	13'h1d85: q3 = 16'h000d; // 0x3b0a
	13'h1d86: q3 = 16'hffeb; // 0x3b0c
	13'h1d87: q3 = 16'hfff5; // 0x3b0e
	13'h1d88: q3 = 16'h0022; // 0x3b10
	13'h1d89: q3 = 16'hffe0; // 0x3b12
	13'h1d8a: q3 = 16'hffe0; // 0x3b14
	13'h1d8b: q3 = 16'h0004; // 0x3b16
	13'h1d8c: q3 = 16'h0000; // 0x3b18
	13'h1d8d: q3 = 16'h0000; // 0x3b1a
	13'h1d8e: q3 = 16'h0000; // 0x3b1c
	13'h1d8f: q3 = 16'h0080; // 0x3b1e
	13'h1d90: q3 = 16'h003a; // 0x3b20
	13'h1d91: q3 = 16'h00e0; // 0x3b22
	13'h1d92: q3 = 16'h0000; // 0x3b24
	13'h1d93: q3 = 16'h0000; // 0x3b26
	13'h1d94: q3 = 16'h8136; // 0x3b28
	13'h1d95: q3 = 16'h0000; // 0x3b2a
	13'h1d96: q3 = 16'hfb00; // 0x3b2c
	13'h1d97: q3 = 16'h0180; // 0x3b2e
	13'h1d98: q3 = 16'h0000; // 0x3b30
	13'h1d99: q3 = 16'h0000; // 0x3b32
	13'h1d9a: q3 = 16'h8136; // 0x3b34
	13'h1d9b: q3 = 16'h0000; // 0x3b36
	13'h1d9c: q3 = 16'hfb06; // 0x3b38
	13'h1d9d: q3 = 16'h0600; // 0x3b3a
	13'h1d9e: q3 = 16'h0000; // 0x3b3c
	13'h1d9f: q3 = 16'h0000; // 0x3b3e
	13'h1da0: q3 = 16'hfb1e; // 0x3b40
	13'h1da1: q3 = 16'h00e0; // 0x3b42
	13'h1da2: q3 = 16'h0000; // 0x3b44
	13'h1da3: q3 = 16'h038e; // 0x3b46
	13'h1da4: q3 = 16'h0000; // 0x3b48
	13'h1da5: q3 = 16'h0000; // 0x3b4a
	13'h1da6: q3 = 16'hfb26; // 0x3b4c
	13'h1da7: q3 = 16'hffff; // 0x3b4e
	13'h1da8: q3 = 16'h0600; // 0x3b50
	13'h1da9: q3 = 16'h0600; // 0x3b52
	13'h1daa: q3 = 16'h0003; // 0x3b54
	13'h1dab: q3 = 16'hf354; // 0x3b56
	13'h1dac: q3 = 16'hf356; // 0x3b58
	13'h1dad: q3 = 16'h0003; // 0x3b5a
	13'h1dae: q3 = 16'h1656; // 0x3b5c
	13'h1daf: q3 = 16'h1655; // 0x3b5e
	13'h1db0: q3 = 16'h0003; // 0x3b60
	13'h1db1: q3 = 16'hcf00; // 0x3b62
	13'h1db2: q3 = 16'hcf00; // 0x3b64
	13'h1db3: q3 = 16'h0001; // 0x3b66
	13'h1db4: q3 = 16'h0a80; // 0x3b68
	13'h1db5: q3 = 16'h0a80; // 0x3b6a
	13'h1db6: q3 = 16'h0004; // 0x3b6c
	13'h1db7: q3 = 16'hec54; // 0x3b6e
	13'h1db8: q3 = 16'hec56; // 0x3b70
	13'h1db9: q3 = 16'h0003; // 0x3b72
	13'h1dba: q3 = 16'h04de; // 0x3b74
	13'h1dbb: q3 = 16'h04db; // 0x3b76
	13'h1dbc: q3 = 16'h0007; // 0x3b78
	13'h1dbd: q3 = 16'hf854; // 0x3b7a
	13'h1dbe: q3 = 16'hf856; // 0x3b7c
	13'h1dbf: q3 = 16'h0003; // 0x3b7e
	13'h1dc0: q3 = 16'h0340; // 0x3b80
	13'h1dc1: q3 = 16'h0340; // 0x3b82
	13'h1dc2: q3 = 16'h0004; // 0x3b84
	13'h1dc3: q3 = 16'hfd60; // 0x3b86
	13'h1dc4: q3 = 16'hfd60; // 0x3b88
	13'h1dc5: q3 = 16'h0008; // 0x3b8a
	13'h1dc6: q3 = 16'h0c56; // 0x3b8c
	13'h1dc7: q3 = 16'h0c55; // 0x3b8e
	13'h1dc8: q3 = 16'h0003; // 0x3b90
	13'h1dc9: q3 = 16'hed00; // 0x3b92
	13'h1dca: q3 = 16'hed00; // 0x3b94
	13'h1dcb: q3 = 16'h0001; // 0x3b96
	13'h1dcc: q3 = 16'h0100; // 0x3b98
	13'h1dcd: q3 = 16'h0100; // 0x3b9a
	13'h1dce: q3 = 16'h0002; // 0x3b9c
	13'h1dcf: q3 = 16'h1500; // 0x3b9e
	13'h1dd0: q3 = 16'h1500; // 0x3ba0
	13'h1dd1: q3 = 16'h0001; // 0x3ba2
	13'h1dd2: q3 = 16'h0100; // 0x3ba4
	13'h1dd3: q3 = 16'h0100; // 0x3ba6
	13'h1dd4: q3 = 16'h0002; // 0x3ba8
	13'h1dd5: q3 = 16'hed00; // 0x3baa
	13'h1dd6: q3 = 16'hed00; // 0x3bac
	13'h1dd7: q3 = 16'h0001; // 0x3bae
	13'h1dd8: q3 = 16'h0356; // 0x3bb0
	13'h1dd9: q3 = 16'h0355; // 0x3bb2
	13'h1dda: q3 = 16'h0003; // 0x3bb4
	13'h1ddb: q3 = 16'heb00; // 0x3bb6
	13'h1ddc: q3 = 16'heb00; // 0x3bb8
	13'h1ddd: q3 = 16'h0001; // 0x3bba
	13'h1dde: q3 = 16'h0456; // 0x3bbc
	13'h1ddf: q3 = 16'h0455; // 0x3bbe
	13'h1de0: q3 = 16'h0003; // 0x3bc0
	13'h1de1: q3 = 16'he200; // 0x3bc2
	13'h1de2: q3 = 16'he200; // 0x3bc4
	13'h1de3: q3 = 16'h0001; // 0x3bc6
	13'h1de4: q3 = 16'h1500; // 0x3bc8
	13'h1de5: q3 = 16'h1500; // 0x3bca
	13'h1de6: q3 = 16'h0001; // 0x3bcc
	13'h1de7: q3 = 16'hf200; // 0x3bce
	13'h1de8: q3 = 16'hf200; // 0x3bd0
	13'h1de9: q3 = 16'h0001; // 0x3bd2
	13'h1dea: q3 = 16'h0180; // 0x3bd4
	13'h1deb: q3 = 16'h0180; // 0x3bd6
	13'h1dec: q3 = 16'h0002; // 0x3bd8
	13'h1ded: q3 = 16'h0480; // 0x3bda
	13'h1dee: q3 = 16'h0480; // 0x3bdc
	13'h1def: q3 = 16'h0002; // 0x3bde
	13'h1df0: q3 = 16'h0380; // 0x3be0
	13'h1df1: q3 = 16'h0380; // 0x3be2
	13'h1df2: q3 = 16'h0004; // 0x3be4
	13'h1df3: q3 = 16'hfa00; // 0x3be6
	13'h1df4: q3 = 16'hfa00; // 0x3be8
	13'h1df5: q3 = 16'h0004; // 0x3bea
	13'h1df6: q3 = 16'h0c00; // 0x3bec
	13'h1df7: q3 = 16'h0c00; // 0x3bee
	13'h1df8: q3 = 16'h0001; // 0x3bf0
	13'h1df9: q3 = 16'h029c; // 0x3bf2
	13'h1dfa: q3 = 16'h0299; // 0x3bf4
	13'h1dfb: q3 = 16'h0005; // 0x3bf6
	13'h1dfc: q3 = 16'hde00; // 0x3bf8
	13'h1dfd: q3 = 16'hde00; // 0x3bfa
	13'h1dfe: q3 = 16'h0001; // 0x3bfc
	13'h1dff: q3 = 16'h0634; // 0x3bfe
	13'h1e00: q3 = 16'h0633; // 0x3c00
	13'h1e01: q3 = 16'h0005; // 0x3c02
	13'h1e02: q3 = 16'he400; // 0x3c04
	13'h1e03: q3 = 16'he400; // 0x3c06
	13'h1e04: q3 = 16'h0001; // 0x3c08
	13'h1e05: q3 = 16'h0b00; // 0x3c0a
	13'h1e06: q3 = 16'h0b00; // 0x3c0c
	13'h1e07: q3 = 16'h0003; // 0x3c0e
	13'h1e08: q3 = 16'hf780; // 0x3c10
	13'h1e09: q3 = 16'hf780; // 0x3c12
	13'h1e0a: q3 = 16'h0002; // 0x3c14
	13'h1e0b: q3 = 16'h0000; // 0x3c16
	13'h1e0c: q3 = 16'h0000; // 0x3c18
	13'h1e0d: q3 = 16'h0000; // 0x3c1a
	13'h1e0e: q3 = 16'h00d8; // 0x3c1c
	13'h1e0f: q3 = 16'h00d5; // 0x3c1e
	13'h1e10: q3 = 16'h0009; // 0x3c20
	13'h1e11: q3 = 16'hffe0; // 0x3c22
	13'h1e12: q3 = 16'hffe0; // 0x3c24
	13'h1e13: q3 = 16'h001c; // 0x3c26
	13'h1e14: q3 = 16'hffc0; // 0x3c28
	13'h1e15: q3 = 16'hffec; // 0x3c2a
	13'h1e16: q3 = 16'h0031; // 0x3c2c
	13'h1e17: q3 = 16'h0000; // 0x3c2e
	13'h1e18: q3 = 16'h0600; // 0x3c30
	13'h1e19: q3 = 16'h0000; // 0x3c32
	13'h1e1a: q3 = 16'h0000; // 0x3c34
	13'h1e1b: q3 = 16'h8136; // 0x3c36
	13'h1e1c: q3 = 16'h0000; // 0x3c38
	13'h1e1d: q3 = 16'hfb50; // 0x3c3a
	13'h1e1e: q3 = 16'h1400; // 0x3c3c
	13'h1e1f: q3 = 16'h0000; // 0x3c3e
	13'h1e20: q3 = 16'h0000; // 0x3c40
	13'h1e21: q3 = 16'h8136; // 0x3c42
	13'h1e22: q3 = 16'h0000; // 0x3c44
	13'h1e23: q3 = 16'hfc1c; // 0x3c46
	13'h1e24: q3 = 16'h0000; // 0x3c48
	13'h1e25: q3 = 16'h0000; // 0x3c4a
	13'h1e26: q3 = 16'h0000; // 0x3c4c
	13'h1e27: q3 = 16'h0000; // 0x3c4e
	13'h1e28: q3 = 16'h00e0; // 0x3c50
	13'h1e29: q3 = 16'h0000; // 0x3c52
	13'h1e2a: q3 = 16'h0514; // 0x3c54
	13'h1e2b: q3 = 16'h0000; // 0x3c56
	13'h1e2c: q3 = 16'h0000; // 0x3c58
	13'h1e2d: q3 = 16'hfc34; // 0x3c5a
	13'h1e2e: q3 = 16'hffff; // 0x3c5c
	13'h1e2f: q3 = 16'h3e00; // 0x3c5e
	13'h1e30: q3 = 16'h362d; // 0x3c60
	13'h1e31: q3 = 16'h3139; // 0x3c62
	13'h1e32: q3 = 16'h362d; // 0x3c64
	13'h1e33: q3 = 16'h3136; // 0x3c66
	13'h1e34: q3 = 16'h2d31; // 0x3c68
	13'h1e35: q3 = 16'h3936; // 0x3c6a
	13'h1e36: q3 = 16'h2d31; // 0x3c6c
	13'h1e37: q3 = 16'h3039; // 0x3c6e
	13'h1e38: q3 = 16'h3136; // 0x3c70
	13'h1e39: q3 = 16'h2d31; // 0x3c72
	13'h1e3a: q3 = 16'h3039; // 0x3c74
	13'h1e3b: q3 = 16'h2d00; // 0x3c76
	13'h1e3c: q3 = 16'h3139; // 0x3c78
	13'h1e3d: q3 = 16'h0000; // 0x3c7a
	13'h1e3e: q3 = 16'hac6e; // 0x3c7c
	13'h1e3f: q3 = 16'h0000; // 0x3c7e
	13'h1e40: q3 = 16'hac66; // 0x3c80
	13'h1e41: q3 = 16'h0000; // 0x3c82
	13'h1e42: q3 = 16'hac8e; // 0x3c84
	13'h1e43: q3 = 16'h0000; // 0x3c86
	13'h1e44: q3 = 16'hac38; // 0x3c88
	13'h1e45: q3 = 16'h0000; // 0x3c8a
	13'h1e46: q3 = 16'hac34; // 0x3c8c
	13'h1e47: q3 = 16'h0000; // 0x3c8e
	13'h1e48: q3 = 16'hac2c; // 0x3c90
	13'h1e49: q3 = 16'h0000; // 0x3c92
	13'h1e4a: q3 = 16'habf4; // 0x3c94
	13'h1e4b: q3 = 16'h0000; // 0x3c96
	13'h1e4c: q3 = 16'habce; // 0x3c98
	13'h1e4d: q3 = 16'h0000; // 0x3c9a
	13'h1e4e: q3 = 16'hac8e; // 0x3c9c
	13'h1e4f: q3 = 16'h0000; // 0x3c9e
	13'h1e50: q3 = 16'hab82; // 0x3ca0
	13'h1e51: q3 = 16'h0000; // 0x3ca2
	13'h1e52: q3 = 16'hab6c; // 0x3ca4
	13'h1e53: q3 = 16'h0000; // 0x3ca6
	13'h1e54: q3 = 16'hab62; // 0x3ca8
	13'h1e55: q3 = 16'h0000; // 0x3caa
	13'h1e56: q3 = 16'hab58; // 0x3cac
	13'h1e57: q3 = 16'h0000; // 0x3cae
	13'h1e58: q3 = 16'hab4e; // 0x3cb0
	13'h1e59: q3 = 16'h0000; // 0x3cb2
	13'h1e5a: q3 = 16'hac8e; // 0x3cb4
	13'h1e5b: q3 = 16'h0000; // 0x3cb6
	13'h1e5c: q3 = 16'hab3e; // 0x3cb8
	13'h1e5d: q3 = 16'h0000; // 0x3cba
	13'h1e5e: q3 = 16'hab34; // 0x3cbc
	13'h1e5f: q3 = 16'h0000; // 0x3cbe
	13'h1e60: q3 = 16'hab2a; // 0x3cc0
	13'h1e61: q3 = 16'h0000; // 0x3cc2
	13'h1e62: q3 = 16'hac8e; // 0x3cc4
	13'h1e63: q3 = 16'h0000; // 0x3cc6
	13'h1e64: q3 = 16'hab20; // 0x3cc8
	13'h1e65: q3 = 16'h0000; // 0x3cca
	13'h1e66: q3 = 16'hab16; // 0x3ccc
	13'h1e67: q3 = 16'h0000; // 0x3cce
	13'h1e68: q3 = 16'hac8e; // 0x3cd0
	13'h1e69: q3 = 16'h0000; // 0x3cd2
	13'h1e6a: q3 = 16'haaf6; // 0x3cd4
	13'h1e6b: q3 = 16'h0000; // 0x3cd6
	13'h1e6c: q3 = 16'haaec; // 0x3cd8
	13'h1e6d: q3 = 16'h0000; // 0x3cda
	13'h1e6e: q3 = 16'haae2; // 0x3cdc
	13'h1e6f: q3 = 16'h2000; // 0x3cde
	13'h1e70: q3 = 16'h2500; // 0x3ce0
	13'h1e71: q3 = 16'h0000; // 0x3ce2
	13'h1e72: q3 = 16'h0000; // 0x3ce4
	13'h1e73: q3 = 16'h0000; // 0x3ce6
	13'h1e74: q3 = 16'hff28; // 0x3ce8
	13'h1e75: q3 = 16'hff2b; // 0x3cea
	13'h1e76: q3 = 16'h0009; // 0x3cec
	13'h1e77: q3 = 16'h0000; // 0x3cee
	13'h1e78: q3 = 16'h0000; // 0x3cf0
	13'h1e79: q3 = 16'h0000; // 0x3cf2
	13'h1e7a: q3 = 16'h00c0; // 0x3cf4
	13'h1e7b: q3 = 16'h0014; // 0x3cf6
	13'h1e7c: q3 = 16'h00e0; // 0x3cf8
	13'h1e7d: q3 = 16'h0000; // 0x3cfa
	13'h1e7e: q3 = 16'h0000; // 0x3cfc
	13'h1e7f: q3 = 16'h8136; // 0x3cfe
	13'h1e80: q3 = 16'h0000; // 0x3d00
	13'h1e81: q3 = 16'hfce2; // 0x3d02
	13'h1e82: q3 = 16'h1800; // 0x3d04
	13'h1e83: q3 = 16'h0000; // 0x3d06
	13'h1e84: q3 = 16'h0000; // 0x3d08
	13'h1e85: q3 = 16'h8136; // 0x3d0a
	13'h1e86: q3 = 16'h0000; // 0x3d0c
	13'h1e87: q3 = 16'hfce8; // 0x3d0e
	13'h1e88: q3 = 16'h0780; // 0x3d10
	13'h1e89: q3 = 16'h0000; // 0x3d12
	13'h1e8a: q3 = 16'h0000; // 0x3d14
	13'h1e8b: q3 = 16'hfcf4; // 0x3d16
	13'h1e8c: q3 = 16'h00e0; // 0x3d18
	13'h1e8d: q3 = 16'h0000; // 0x3d1a
	13'h1e8e: q3 = 16'h05aa; // 0x3d1c
	13'h1e8f: q3 = 16'h0000; // 0x3d1e
	13'h1e90: q3 = 16'h0000; // 0x3d20
	13'h1e91: q3 = 16'hfcfc; // 0x3d22
	13'h1e92: q3 = 16'hffff; // 0x3d24
	13'h1e93: q3 = 16'h0000; // 0x3d26
	13'h1e94: q3 = 16'hb2d6; // 0x3d28
	13'h1e95: q3 = 16'h0000; // 0x3d2a
	13'h1e96: q3 = 16'hb2e4; // 0x3d2c
	13'h1e97: q3 = 16'h0000; // 0x3d2e
	13'h1e98: q3 = 16'hb2f0; // 0x3d30
	13'h1e99: q3 = 16'h0000; // 0x3d32
	13'h1e9a: q3 = 16'hb2fe; // 0x3d34
	13'h1e9b: q3 = 16'h0000; // 0x3d36
	13'h1e9c: q3 = 16'hb30c; // 0x3d38
	13'h1e9d: q3 = 16'h0000; // 0x3d3a
	13'h1e9e: q3 = 16'hb314; // 0x3d3c
	13'h1e9f: q3 = 16'h0000; // 0x3d3e
	13'h1ea0: q3 = 16'hb31c; // 0x3d40
	13'h1ea1: q3 = 16'h0000; // 0x3d42
	13'h1ea2: q3 = 16'hb324; // 0x3d44
	13'h1ea3: q3 = 16'h0000; // 0x3d46
	13'h1ea4: q3 = 16'hb32c; // 0x3d48
	13'h1ea5: q3 = 16'h0000; // 0x3d4a
	13'h1ea6: q3 = 16'hb334; // 0x3d4c
	13'h1ea7: q3 = 16'hfde0; // 0x3d4e
	13'h1ea8: q3 = 16'hfde0; // 0x3d50
	13'h1ea9: q3 = 16'h003c; // 0x3d52
	13'h1eaa: q3 = 16'h0000; // 0x3d54
	13'h1eab: q3 = 16'h0000; // 0x3d56
	13'h1eac: q3 = 16'h0000; // 0x3d58
	13'h1ead: q3 = 16'h0080; // 0x3d5a
	13'h1eae: q3 = 16'h0080; // 0x3d5c
	13'h1eaf: q3 = 16'h000f; // 0x3d5e
	13'h1eb0: q3 = 16'h0000; // 0x3d60
	13'h1eb1: q3 = 16'h0000; // 0x3d62
	13'h1eb2: q3 = 16'h002c; // 0x3d64
	13'h1eb3: q3 = 16'hf880; // 0x3d66
	13'h1eb4: q3 = 16'hf880; // 0x3d68
	13'h1eb5: q3 = 16'h0001; // 0x3d6a
	13'h1eb6: q3 = 16'h0000; // 0x3d6c
	13'h1eb7: q3 = 16'h0000; // 0x3d6e
	13'h1eb8: q3 = 16'h7fff; // 0x3d70
	13'h1eb9: q3 = 16'h0000; // 0x3d72
	13'h1eba: q3 = 16'h8136; // 0x3d74
	13'h1ebb: q3 = 16'h0000; // 0x3d76
	13'h1ebc: q3 = 16'hfd4e; // 0x3d78
	13'h1ebd: q3 = 16'h7f80; // 0x3d7a
	13'h1ebe: q3 = 16'h0000; // 0x3d7c
	13'h1ebf: q3 = 16'h0000; // 0x3d7e
	13'h1ec0: q3 = 16'h8136; // 0x3d80
	13'h1ec1: q3 = 16'h0000; // 0x3d82
	13'h1ec2: q3 = 16'hfd5a; // 0x3d84
	13'h1ec3: q3 = 16'h0000; // 0x3d86
	13'h1ec4: q3 = 16'h0000; // 0x3d88
	13'h1ec5: q3 = 16'h0000; // 0x3d8a
	13'h1ec6: q3 = 16'h0000; // 0x3d8c
	13'h1ec7: q3 = 16'h00e0; // 0x3d8e
	13'h1ec8: q3 = 16'h0000; // 0x3d90
	13'h1ec9: q3 = 16'h1388; // 0x3d92
	13'h1eca: q3 = 16'h0000; // 0x3d94
	13'h1ecb: q3 = 16'h0000; // 0x3d96
	13'h1ecc: q3 = 16'hfd72; // 0x3d98
	13'h1ecd: q3 = 16'hffff; // 0x3d9a
	13'h1ece: q3 = 16'hfdda; // 0x3d9c
	13'h1ecf: q3 = 16'hfde3; // 0x3d9e
	13'h1ed0: q3 = 16'h0023; // 0x3da0
	13'h1ed1: q3 = 16'h00cf; // 0x3da2
	13'h1ed2: q3 = 16'h00c9; // 0x3da4
	13'h1ed3: q3 = 16'h002a; // 0x3da6
	13'h1ed4: q3 = 16'h0000; // 0x3da8
	13'h1ed5: q3 = 16'h0000; // 0x3daa
	13'h1ed6: q3 = 16'h0000; // 0x3dac
	13'h1ed7: q3 = 16'h0038; // 0x3dae
	13'h1ed8: q3 = 16'h0018; // 0x3db0
	13'h1ed9: q3 = 16'h0024; // 0x3db2
	13'h1eda: q3 = 16'hffda; // 0x3db4
	13'h1edb: q3 = 16'hffea; // 0x3db6
	13'h1edc: q3 = 16'h0028; // 0x3db8
	13'h1edd: q3 = 16'h0000; // 0x3dba
	13'h1ede: q3 = 16'hfdda; // 0x3dbc
	13'h1edf: q3 = 16'h0000; // 0x3dbe
	13'h1ee0: q3 = 16'h0080; // 0x3dc0
	13'h1ee1: q3 = 16'h0059; // 0x3dc2
	13'h1ee2: q3 = 16'h00e0; // 0x3dc4
	13'h1ee3: q3 = 16'h0000; // 0x3dc6
	13'h1ee4: q3 = 16'h0000; // 0x3dc8
	13'h1ee5: q3 = 16'h8136; // 0x3dca
	13'h1ee6: q3 = 16'h0000; // 0x3dcc
	13'h1ee7: q3 = 16'hfd9c; // 0x3dce
	13'h1ee8: q3 = 16'h5b00; // 0x3dd0
	13'h1ee9: q3 = 16'h0000; // 0x3dd2
	13'h1eea: q3 = 16'h0000; // 0x3dd4
	13'h1eeb: q3 = 16'h8136; // 0x3dd6
	13'h1eec: q3 = 16'h0000; // 0x3dd8
	13'h1eed: q3 = 16'hfdae; // 0x3dda
	13'h1eee: q3 = 16'h0000; // 0x3ddc
	13'h1eef: q3 = 16'h0000; // 0x3dde
	13'h1ef0: q3 = 16'h0000; // 0x3de0
	13'h1ef1: q3 = 16'hfdc0; // 0x3de2
	13'h1ef2: q3 = 16'h00e0; // 0x3de4
	13'h1ef3: q3 = 16'h0000; // 0x3de6
	13'h1ef4: q3 = 16'h0040; // 0x3de8
	13'h1ef5: q3 = 16'h0058; // 0x3dea
	13'h1ef6: q3 = 16'h0000; // 0x3dec
	13'h1ef7: q3 = 16'h0000; // 0x3dee
	13'h1ef8: q3 = 16'h0000; // 0x3df0
	13'h1ef9: q3 = 16'hfde8; // 0x3df2
	13'h1efa: q3 = 16'h0000; // 0x3df4
	13'h1efb: q3 = 16'h0000; // 0x3df6
	13'h1efc: q3 = 16'h0578; // 0x3df8
	13'h1efd: q3 = 16'h0001; // 0x3dfa
	13'h1efe: q3 = 16'h0000; // 0x3dfc
	13'h1eff: q3 = 16'hfdc8; // 0x3dfe
	13'h1f00: q3 = 16'h0000; // 0x3e00
	13'h1f01: q3 = 16'hfdf0; // 0x3e02
	13'h1f02: q3 = 16'hffff; // 0x3e04
	13'h1f03: q3 = 16'h0808; // 0x3e06
	13'h1f04: q3 = 16'h0800; // 0x3e08
	13'h1f05: q3 = 16'h0000; // 0x3e0a
	13'h1f06: q3 = 16'h0000; // 0x3e0c
	13'h1f07: q3 = 16'h0011; // 0x3e0e
	13'h1f08: q3 = 16'h1111; // 0x3e10
	13'h1f09: q3 = 16'h1111; // 0x3e12
	13'h1f0a: q3 = 16'h1100; // 0x3e14
	13'h1f0b: q3 = 16'h1513; // 0x3e16
	13'h1f0c: q3 = 16'h110f; // 0x3e18
	13'h1f0d: q3 = 16'h0d0b; // 0x3e1a
	13'h1f0e: q3 = 16'h0907; // 0x3e1c
	13'h1f0f: q3 = 16'h050f; // 0x3e1e
	13'h1f10: q3 = 16'h0d0b; // 0x3e20
	13'h1f11: q3 = 16'h0907; // 0x3e22
	13'h1f12: q3 = 16'h0500; // 0x3e24
	13'h1f13: q3 = 16'h4641; // 0x3e26
	13'h1f14: q3 = 16'h4255; // 0x3e28
	13'h1f15: q3 = 16'h4c4f; // 0x3e2a
	13'h1f16: q3 = 16'h5553; // 0x3e2c
	13'h1f17: q3 = 16'h2046; // 0x3e2e
	13'h1f18: q3 = 16'h4f4f; // 0x3e30
	13'h1f19: q3 = 16'h4420; // 0x3e32
	13'h1f1a: q3 = 16'h464c; // 0x3e34
	13'h1f1b: q3 = 16'h494e; // 0x3e36
	13'h1f1c: q3 = 16'h4745; // 0x3e38
	13'h1f1d: q3 = 16'h5253; // 0x3e3a
	13'h1f1e: q3 = 16'h0020; // 0x3e3c
	13'h1f1f: q3 = 16'h0020; // 0x3e3e
	13'h1f20: q3 = 16'h0030; // 0x3e40
	13'h1f21: q3 = 16'h3000; // 0x3e42
	13'h1f22: q3 = 16'h0000; // 0x3e44
	13'h1f23: q3 = 16'h003c; // 0x3e46
	13'h1f24: q3 = 16'h3000; // 0x3e48
	13'h1f25: q3 = 16'h3030; // 0x3e4a
	13'h1f26: q3 = 16'h003a; // 0x3e4c
	13'h1f27: q3 = 16'h0000; // 0x3e4e
	13'h1f28: q3 = 16'h0000; // 0x3e50
	13'h1f29: q3 = 16'hbb1e; // 0x3e52
	13'h1f2a: q3 = 16'h0000; // 0x3e54
	13'h1f2b: q3 = 16'hbb96; // 0x3e56
	13'h1f2c: q3 = 16'h0000; // 0x3e58
	13'h1f2d: q3 = 16'hbbac; // 0x3e5a
	13'h1f2e: q3 = 16'h0000; // 0x3e5c
	13'h1f2f: q3 = 16'hbbc0; // 0x3e5e
	13'h1f30: q3 = 16'h0000; // 0x3e60
	13'h1f31: q3 = 16'hbbdc; // 0x3e62
	13'h1f32: q3 = 16'h0000; // 0x3e64
	13'h1f33: q3 = 16'hbbe0; // 0x3e66
	13'h1f34: q3 = 16'h0000; // 0x3e68
	13'h1f35: q3 = 16'hbbe4; // 0x3e6a
	13'h1f36: q3 = 16'h0000; // 0x3e6c
	13'h1f37: q3 = 16'hbc0e; // 0x3e6e
	13'h1f38: q3 = 16'h0000; // 0x3e70
	13'h1f39: q3 = 16'hbcf6; // 0x3e72
	13'h1f3a: q3 = 16'h0000; // 0x3e74
	13'h1f3b: q3 = 16'hbd14; // 0x3e76
	13'h1f3c: q3 = 16'h0000; // 0x3e78
	13'h1f3d: q3 = 16'hbd2a; // 0x3e7a
	13'h1f3e: q3 = 16'h0000; // 0x3e7c
	13'h1f3f: q3 = 16'hbd3c; // 0x3e7e
	13'h1f40: q3 = 16'h0000; // 0x3e80
	13'h1f41: q3 = 16'hbd46; // 0x3e82
	13'h1f42: q3 = 16'h0000; // 0x3e84
	13'h1f43: q3 = 16'hbd50; // 0x3e86
	13'h1f44: q3 = 16'h0000; // 0x3e88
	13'h1f45: q3 = 16'hbd7e; // 0x3e8a
	13'h1f46: q3 = 16'h0000; // 0x3e8c
	13'h1f47: q3 = 16'hbd98; // 0x3e8e
	13'h1f48: q3 = 16'h005a; // 0x3e90
	13'h1f49: q3 = 16'h004b; // 0x3e92
	13'h1f4a: q3 = 16'h0033; // 0x3e94
	13'h1f4b: q3 = 16'h00d0; // 0x3e96
	13'h1f4c: q3 = 16'h00ac; // 0x3e98
	13'h1f4d: q3 = 16'h0025; // 0x3e9a
	13'h1f4e: q3 = 16'h0000; // 0x3e9c
	13'h1f4f: q3 = 16'h0000; // 0x3e9e
	13'h1f50: q3 = 16'h0000; // 0x3ea0
	13'h1f51: q3 = 16'h0140; // 0x3ea2
	13'h1f52: q3 = 16'h0140; // 0x3ea4
	13'h1f53: q3 = 16'h0006; // 0x3ea6
	13'h1f54: q3 = 16'hffc7; // 0x3ea8
	13'h1f55: q3 = 16'hffe9; // 0x3eaa
	13'h1f56: q3 = 16'h0052; // 0x3eac
	13'h1f57: q3 = 16'h0000; // 0x3eae
	13'h1f58: q3 = 16'h005a; // 0x3eb0
	13'h1f59: q3 = 16'h0000; // 0x3eb2
	13'h1f5a: q3 = 16'h0000; // 0x3eb4
	13'h1f5b: q3 = 16'h8136; // 0x3eb6
	13'h1f5c: q3 = 16'h0000; // 0x3eb8
	13'h1f5d: q3 = 16'hfe90; // 0x3eba
	13'h1f5e: q3 = 16'h0900; // 0x3ebc
	13'h1f5f: q3 = 16'h0000; // 0x3ebe
	13'h1f60: q3 = 16'h0000; // 0x3ec0
	13'h1f61: q3 = 16'h8136; // 0x3ec2
	13'h1f62: q3 = 16'h0000; // 0x3ec4
	13'h1f63: q3 = 16'hfea2; // 0x3ec6
	13'h1f64: q3 = 16'h0000; // 0x3ec8
	13'h1f65: q3 = 16'h0000; // 0x3eca
	13'h1f66: q3 = 16'h0000; // 0x3ecc
	13'h1f67: q3 = 16'h0000; // 0x3ece
	13'h1f68: q3 = 16'h00e0; // 0x3ed0
	13'h1f69: q3 = 16'h0000; // 0x3ed2
	13'h1f6a: q3 = 16'h05d2; // 0x3ed4
	13'h1f6b: q3 = 16'h0000; // 0x3ed6
	13'h1f6c: q3 = 16'h0000; // 0x3ed8
	13'h1f6d: q3 = 16'hfeb4; // 0x3eda
	13'h1f6e: q3 = 16'hffff; // 0x3edc
	13'h1f6f: q3 = 16'hff86; // 0x3ede
	13'h1f70: q3 = 16'hffaa; // 0x3ee0
	13'h1f71: q3 = 16'h004a; // 0x3ee2
	13'h1f72: q3 = 16'hff99; // 0x3ee4
	13'h1f73: q3 = 16'hffdb; // 0x3ee6
	13'h1f74: q3 = 16'h0066; // 0x3ee8
	13'h1f75: q3 = 16'h0000; // 0x3eea
	13'h1f76: q3 = 16'h0000; // 0x3eec
	13'h1f77: q3 = 16'h0000; // 0x3eee
	13'h1f78: q3 = 16'h003c; // 0x3ef0
	13'h1f79: q3 = 16'h0009; // 0x3ef2
	13'h1f7a: q3 = 16'h00a5; // 0x3ef4
	13'h1f7b: q3 = 16'hff4c; // 0x3ef6
	13'h1f7c: q3 = 16'hff52; // 0x3ef8
	13'h1f7d: q3 = 16'h000b; // 0x3efa
	13'h1f7e: q3 = 16'h0000; // 0x3efc
	13'h1f7f: q3 = 16'hff86; // 0x3efe
	13'h1f80: q3 = 16'h0000; // 0x3f00
	13'h1f81: q3 = 16'h0000; // 0x3f02
	13'h1f82: q3 = 16'h8136; // 0x3f04
	13'h1f83: q3 = 16'h0000; // 0x3f06
	13'h1f84: q3 = 16'hfede; // 0x3f08
	13'h1f85: q3 = 16'h3100; // 0x3f0a
	13'h1f86: q3 = 16'h0000; // 0x3f0c
	13'h1f87: q3 = 16'h0000; // 0x3f0e
	13'h1f88: q3 = 16'h8136; // 0x3f10
	13'h1f89: q3 = 16'h0000; // 0x3f12
	13'h1f8a: q3 = 16'hfef0; // 0x3f14
	13'h1f8b: q3 = 16'h0180; // 0x3f16
	13'h1f8c: q3 = 16'h0000; // 0x3f18
	13'h1f8d: q3 = 16'h0000; // 0x3f1a
	13'h1f8e: q3 = 16'h0000; // 0x3f1c
	13'h1f8f: q3 = 16'h00e0; // 0x3f1e
	13'h1f90: q3 = 16'h0000; // 0x3f20
	13'h1f91: q3 = 16'h05dc; // 0x3f22
	13'h1f92: q3 = 16'h0000; // 0x3f24
	13'h1f93: q3 = 16'h0000; // 0x3f26
	13'h1f94: q3 = 16'hff02; // 0x3f28
	13'h1f95: q3 = 16'hffff; // 0x3f2a
	13'h1f96: q3 = 16'h46fc; // 0x3f2c
	13'h1f97: q3 = 16'h2700; // 0x3f2e
	13'h1f98: q3 = 16'h4a79; // 0x3f30
	13'h1f99: q3 = 16'h0095; // 0x3f32
	13'h1f9a: q3 = 16'h8000; // 0x3f34
	13'h1f9b: q3 = 16'h2e79; // 0x3f36
	13'h1f9c: q3 = 16'h0000; // 0x3f38
	13'h1f9d: q3 = 16'h0000; // 0x3f3a
	13'h1f9e: q3 = 16'h227c; // 0x3f3c
	13'h1f9f: q3 = 16'h0000; // 0x3f3e
	13'h1fa0: q3 = 16'h04e0; // 0x3f40
	13'h1fa1: q3 = 16'h247c; // 0x3f42
	13'h1fa2: q3 = 16'h0000; // 0x3f44
	13'h1fa3: q3 = 16'h04e8; // 0x3f46
	13'h1fa4: q3 = 16'h4a79; // 0x3f48
	13'h1fa5: q3 = 16'h0095; // 0x3f4a
	13'h1fa6: q3 = 16'h8000; // 0x3f4c
	13'h1fa7: q3 = 16'hb5c9; // 0x3f4e
	13'h1fa8: q3 = 16'h6d00; // 0x3f50
	13'h1fa9: q3 = 16'h0006; // 0x3f52
	13'h1faa: q3 = 16'h4259; // 0x3f54
	13'h1fab: q3 = 16'h60f0; // 0x3f56
	13'h1fac: q3 = 16'h227c; // 0x3f58
	13'h1fad: q3 = 16'h0000; // 0x3f5a
	13'h1fae: q3 = 16'h04e0; // 0x3f5c
	13'h1faf: q3 = 16'h4281; // 0x3f5e
	13'h1fb0: q3 = 16'h4a79; // 0x3f60
	13'h1fb1: q3 = 16'h0095; // 0x3f62
	13'h1fb2: q3 = 16'h8000; // 0x3f64
	13'h1fb3: q3 = 16'hb279; // 0x3f66
	13'h1fb4: q3 = 16'h0000; // 0x3f68
	13'h1fb5: q3 = 16'h04d6; // 0x3f6a
	13'h1fb6: q3 = 16'h6c00; // 0x3f6c
	13'h1fb7: q3 = 16'h005e; // 0x3f6e
	13'h1fb8: q3 = 16'h2a01; // 0x3f70
	13'h1fb9: q3 = 16'he345; // 0x3f72
	13'h1fba: q3 = 16'he345; // 0x3f74
	13'h1fbb: q3 = 16'h2a7c; // 0x3f76
	13'h1fbc: q3 = 16'h0000; // 0x3f78
	13'h1fbd: q3 = 16'h04dc; // 0x3f7a
	13'h1fbe: q3 = 16'hdbc5; // 0x3f7c
	13'h1fbf: q3 = 16'h2455; // 0x3f7e
	13'h1fc0: q3 = 16'he245; // 0x3f80
	13'h1fc1: q3 = 16'h4242; // 0x3f82
	13'h1fc2: q3 = 16'h4a79; // 0x3f84
	13'h1fc3: q3 = 16'h0095; // 0x3f86
	13'h1fc4: q3 = 16'h8000; // 0x3f88
	13'h1fc5: q3 = 16'h2a7c; // 0x3f8a
	13'h1fc6: q3 = 16'h0000; // 0x3f8c
	13'h1fc7: q3 = 16'h04da; // 0x3f8e
	13'h1fc8: q3 = 16'hdbc5; // 0x3f90
	13'h1fc9: q3 = 16'hb455; // 0x3f92
	13'h1fca: q3 = 16'h6c00; // 0x3f94
	13'h1fcb: q3 = 16'h0032; // 0x3f96
	13'h1fcc: q3 = 16'h4203; // 0x3f98
	13'h1fcd: q3 = 16'h4204; // 0x3f9a
	13'h1fce: q3 = 16'h264a; // 0x3f9c
	13'h1fcf: q3 = 16'h2a7c; // 0x3f9e
	13'h1fd0: q3 = 16'h0000; // 0x3fa0
	13'h1fd1: q3 = 16'h04d8; // 0x3fa2
	13'h1fd2: q3 = 16'hdbc5; // 0x3fa4
	13'h1fd3: q3 = 16'h3c15; // 0x3fa6
	13'h1fd4: q3 = 16'h48c6; // 0x3fa8
	13'h1fd5: q3 = 16'hd7c6; // 0x3faa
	13'h1fd6: q3 = 16'h4246; // 0x3fac
	13'h1fd7: q3 = 16'h4a79; // 0x3fae
	13'h1fd8: q3 = 16'h0095; // 0x3fb0
	13'h1fd9: q3 = 16'h8000; // 0x3fb2
	13'h1fda: q3 = 16'hb5cb; // 0x3fb4
	13'h1fdb: q3 = 16'h6c00; // 0x3fb6
	13'h1fdc: q3 = 16'h0008; // 0x3fb8
	13'h1fdd: q3 = 16'hd61a; // 0x3fba
	13'h1fde: q3 = 16'hd81a; // 0x3fbc
	13'h1fdf: q3 = 16'h60ee; // 0x3fbe
	13'h1fe0: q3 = 16'h12c3; // 0x3fc0
	13'h1fe1: q3 = 16'h12c4; // 0x3fc2
	13'h1fe2: q3 = 16'h5242; // 0x3fc4
	13'h1fe3: q3 = 16'h60bc; // 0x3fc6
	13'h1fe4: q3 = 16'h5241; // 0x3fc8
	13'h1fe5: q3 = 16'h6094; // 0x3fca
	13'h1fe6: q3 = 16'h4241; // 0x3fcc
	13'h1fe7: q3 = 16'h4242; // 0x3fce
	13'h1fe8: q3 = 16'h227c; // 0x3fd0
	13'h1fe9: q3 = 16'h0000; // 0x3fd2
	13'h1fea: q3 = 16'h04e0; // 0x3fd4
	13'h1feb: q3 = 16'h247c; // 0x3fd6
	13'h1fec: q3 = 16'h0000; // 0x3fd8
	13'h1fed: q3 = 16'h04e8; // 0x3fda
	13'h1fee: q3 = 16'h4a79; // 0x3fdc
	13'h1fef: q3 = 16'h0095; // 0x3fde
	13'h1ff0: q3 = 16'h8000; // 0x3fe0
	13'h1ff1: q3 = 16'hb3ca; // 0x3fe2
	13'h1ff2: q3 = 16'h6c00; // 0x3fe4
	13'h1ff3: q3 = 16'h0008; // 0x3fe6
	13'h1ff4: q3 = 16'hd219; // 0x3fe8
	13'h1ff5: q3 = 16'hd419; // 0x3fea
	13'h1ff6: q3 = 16'h60ee; // 0x3fec
	13'h1ff7: q3 = 16'h4401; // 0x3fee
	13'h1ff8: q3 = 16'h4402; // 0x3ff0
	13'h1ff9: q3 = 16'h13c1; // 0x3ff2
	13'h1ffa: q3 = 16'h0000; // 0x3ff4
	13'h1ffb: q3 = 16'h04e8; // 0x3ff6
	13'h1ffc: q3 = 16'h13c2; // 0x3ff8
	13'h1ffd: q3 = 16'h0000; // 0x3ffa
	13'h1ffe: q3 = 16'h04e9; // 0x3ffc
	13'h1fff: q3 = 16'h4ef9; // 0x3ffe
  endcase

  assign out = ~ce0 ? q0 :
               ~ce1 ? q1 :
               ~ce2 ? q2 :
               ~ce3 ? q3 :
               16'h0;

