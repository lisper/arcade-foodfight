    Mac OS X            	   2   �      �                                      ATTR       �   �   F                  �   F  com.apple.quarantine q/0001;53888be4;Google\x20Chrome;1BFB4208-57D9-45D6-956B-B3239B439061 